magic
tech sky130A
magscale 1 2
timestamp 1770726631
<< viali >>
rect 1650 -38 1750 20
rect 3180 -40 3286 10
rect 1662 -1902 1754 -1854
rect 3188 -1908 3280 -1854
<< metal1 >>
rect 3226 712 3490 714
rect 582 408 4394 712
rect 1103 404 1357 408
rect 1146 0 1357 404
rect 1600 20 1800 408
rect 1146 -230 1358 0
rect 1600 -38 1650 20
rect 1750 -38 1800 20
rect 1600 -44 1800 -38
rect 3132 406 3488 408
rect 3132 10 3332 406
rect 3132 -40 3180 10
rect 3286 -40 3332 10
rect 3132 -48 3332 -40
rect 1666 -142 2018 -90
rect 2070 -142 2076 -90
rect 3200 -144 3608 -96
rect 1146 -432 1680 -230
rect 1722 -432 3210 -236
rect 3246 -456 3252 -200
rect 3432 -456 3438 -200
rect 1666 -564 2018 -512
rect 2070 -564 2076 -512
rect 3560 -526 3608 -144
rect 396 -768 596 -700
rect 2018 -768 2070 -564
rect 3202 -574 3608 -526
rect 4329 -565 4414 -561
rect 4796 -565 4996 -524
rect 396 -779 2070 -768
rect 396 -832 2071 -779
rect 396 -842 2070 -832
rect 396 -900 596 -842
rect 400 -1236 600 -1172
rect 400 -1308 1548 -1236
rect 1620 -1308 1626 -1236
rect 400 -1372 600 -1308
rect 2018 -1490 2070 -842
rect 3560 -1236 3608 -574
rect 4328 -567 4996 -565
rect 4328 -652 4329 -567
rect 4414 -652 4996 -567
rect 4329 -658 4414 -652
rect 4796 -724 4996 -652
rect 2108 -1308 2114 -1236
rect 2186 -1308 3608 -1236
rect 1674 -1542 2072 -1490
rect 3560 -1496 3608 -1308
rect 3198 -1536 3608 -1496
rect 3198 -1542 3603 -1536
rect 1217 -1700 1686 -1590
rect 1726 -1607 1798 -1590
rect 1726 -1680 1909 -1607
rect 1982 -1680 1988 -1607
rect 1726 -1698 1798 -1680
rect 1217 -2304 1327 -1700
rect 2020 -1748 2072 -1542
rect 1674 -1800 2072 -1748
rect 2702 -1708 3212 -1604
rect 3434 -1622 3519 -1617
rect 3253 -1623 3519 -1622
rect 3253 -1708 3434 -1623
rect 1620 -1854 1794 -1838
rect 1620 -1902 1662 -1854
rect 1754 -1902 1794 -1854
rect 1620 -2304 1794 -1902
rect 2702 -2304 2806 -1708
rect 3434 -1714 3519 -1708
rect 3557 -1753 3603 -1542
rect 3199 -1799 3603 -1753
rect 3144 -1854 3318 -1848
rect 3144 -1908 3188 -1854
rect 3280 -1908 3318 -1854
rect 3144 -2304 3318 -1908
rect 538 -2608 4350 -2304
<< via1 >>
rect 2018 -142 2070 -90
rect 3252 -456 3432 -200
rect 2018 -564 2070 -512
rect 1548 -1308 1620 -1236
rect 4329 -652 4414 -567
rect 2114 -1308 2186 -1236
rect 1909 -1680 1982 -1607
rect 3434 -1708 3519 -1623
<< metal2 >>
rect 2018 -90 2070 -84
rect 2018 -512 2070 -142
rect 3252 -200 3432 -194
rect 3432 -370 4098 -285
rect 3252 -462 3432 -456
rect 2018 -570 2070 -564
rect 4013 -567 4098 -370
rect 4013 -652 4329 -567
rect 4414 -652 4420 -567
rect 4013 -1010 4098 -652
rect 2333 -1083 4098 -1010
rect 1548 -1236 1620 -1230
rect 2114 -1236 2186 -1230
rect 1620 -1308 2114 -1236
rect 1548 -1314 1620 -1308
rect 2114 -1314 2186 -1308
rect 1909 -1607 1982 -1601
rect 2333 -1607 2406 -1083
rect 1982 -1680 2406 -1607
rect 4013 -1623 4098 -1083
rect 1909 -1686 1982 -1680
rect 3428 -1708 3434 -1623
rect 3519 -1708 4098 -1623
rect 4013 -1718 4098 -1708
use sky130_fd_pr__pfet_01v8_XJP3BL  XM1
timestamp 1770726631
transform 1 0 1701 0 1 -327
box -211 -369 211 369
use sky130_fd_pr__pfet_01v8_XJP3BL  XM2
timestamp 1770726631
transform 1 0 3233 0 1 -333
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_CSX3TK  XM3
timestamp 1770726631
transform 1 0 1707 0 1 -1645
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_CSX3TK  XM4
timestamp 1770726631
transform 1 0 3233 0 1 -1649
box -211 -285 211 285
<< labels >>
flabel metal1 4796 -724 4996 -524 0 FreeSans 256 0 0 0 y
port 2 nsew
flabel metal1 792 490 992 690 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 792 -2572 992 -2372 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 396 -900 596 -700 0 FreeSans 256 0 0 0 a
port 1 nsew
flabel metal1 400 -1372 600 -1172 0 FreeSans 256 0 0 0 b
port 3 nsew
<< end >>
