magic
tech sky130A
magscale 1 2
timestamp 1770730625
<< metal1 >>
rect 874 -1964 2190 -1677
rect 874 -1989 2760 -1964
rect 5974 -1986 8360 -1678
rect 11986 -1991 12821 -1679
rect 6400 -2918 6961 -2916
rect 6400 -2934 7144 -2918
rect 8000 -2934 8200 -2915
rect 1252 -3092 1452 -3090
rect 1252 -3290 2200 -3092
rect 6400 -3095 8200 -2934
rect 6400 -3106 7146 -3095
rect 6400 -3116 7144 -3106
rect 6944 -3118 7144 -3116
rect 1391 -3292 2200 -3290
rect 8000 -3292 8200 -3095
rect 12464 -3535 12563 -3115
rect 1375 -3565 2204 -3564
rect 7535 -3565 8204 -3564
rect 1252 -3764 2204 -3565
rect 7436 -3764 8204 -3565
rect 12458 -3634 12464 -3535
rect 12563 -3634 12569 -3535
rect 1252 -3765 1452 -3764
rect 7436 -3765 7636 -3764
rect 1303 -4458 1402 -3765
rect 1303 -4557 2323 -4458
rect 2422 -4557 2428 -4458
rect 862 -4999 2273 -4696
rect 5501 -4945 5701 -4745
rect 5943 -5005 8156 -4699
rect 11943 -5001 12778 -4689
<< via1 >>
rect 12464 -3634 12563 -3535
rect 2323 -4557 2422 -4458
<< metal2 >>
rect 12464 -3535 12563 -3529
rect 2323 -4458 2422 -4452
rect 12464 -4458 12563 -3634
rect 2422 -4557 12563 -4458
rect 2323 -4563 2422 -4557
use nor_gate  x1
timestamp 1770726631
transform 1 0 1604 0 1 -2392
box 396 -2608 4996 714
use nor_gate  x2
timestamp 1770726631
transform 1 0 7604 0 1 -2392
box 396 -2608 4996 714
<< labels >>
flabel metal1 6386 -1953 6586 -1753 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1252 -3290 1452 -3090 0 FreeSans 256 0 0 0 s
port 1 nsew
flabel metal1 5501 -4945 5701 -4745 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 6944 -3118 7144 -2918 0 FreeSans 256 0 0 0 q
port 3 nsew
flabel metal1 1252 -3765 1452 -3565 0 FreeSans 256 0 0 0 qb
port 2 nsew
flabel metal1 7436 -3765 7636 -3565 0 FreeSans 256 0 0 0 r
port 5 nsew
<< end >>
