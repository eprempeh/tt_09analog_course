magic
tech sky130A
magscale 1 2
timestamp 1771589982
<< metal1 >>
rect 8690 40436 8696 40748
rect 9008 40436 19258 40748
rect 24970 40096 25170 40102
rect 19278 40066 19478 40072
rect 18252 39976 18452 39982
rect 18252 38860 18452 39776
rect 19278 39135 19478 39866
rect 24970 39307 25170 39896
rect 25462 39102 25662 39108
rect 18252 38660 19478 38860
rect 25462 38660 25662 38902
rect 8651 37426 8657 37729
rect 8960 37426 19762 37729
<< via1 >>
rect 8696 40436 9008 40748
rect 18252 39776 18452 39976
rect 19278 39866 19478 40066
rect 24970 39896 25170 40096
rect 25462 38902 25662 39102
rect 8657 37426 8960 37729
<< metal2 >>
rect 18252 42694 18452 42703
rect 8696 40748 9008 40754
rect 5263 40436 5272 40748
rect 5584 40436 8696 40748
rect 8696 40430 9008 40436
rect 18252 39976 18452 42494
rect 19278 42534 27038 42734
rect 27238 42534 27247 42734
rect 19278 40066 19478 42534
rect 25462 42004 25662 42013
rect 23299 41756 23308 41956
rect 23508 41756 25170 41956
rect 24970 40096 25170 41756
rect 18246 39776 18252 39976
rect 18452 39776 18458 39976
rect 19272 39866 19278 40066
rect 19478 39866 19484 40066
rect 24964 39896 24970 40096
rect 25170 39896 25176 40096
rect 25462 39102 25662 41804
rect 25456 38902 25462 39102
rect 25662 38902 25668 39102
rect 8657 37729 8960 37735
rect 5336 37426 5345 37729
rect 5648 37426 8657 37729
rect 8657 37420 8960 37426
<< via2 >>
rect 18252 42494 18452 42694
rect 5272 40436 5584 40748
rect 27038 42534 27238 42734
rect 23308 41756 23508 41956
rect 25462 41804 25662 42004
rect 5345 37426 5648 37729
<< metal3 >>
rect 23306 44116 23506 44122
rect 18252 43508 18452 43514
rect 18252 42699 18452 43308
rect 18247 42694 18457 42699
rect 18247 42494 18252 42694
rect 18452 42494 18457 42694
rect 18247 42489 18457 42494
rect 23306 42162 23506 43916
rect 27038 43190 27238 43196
rect 27038 42739 27238 42990
rect 27033 42734 27243 42739
rect 27033 42534 27038 42734
rect 27238 42534 27243 42734
rect 27033 42529 27243 42534
rect 23306 42090 23508 42162
rect 23308 41961 23508 42090
rect 25457 42004 25667 42009
rect 23303 41956 23513 41961
rect 23303 41756 23308 41956
rect 23508 41756 23513 41956
rect 25457 41804 25462 42004
rect 25662 41804 27580 42004
rect 27780 41804 27786 42004
rect 25457 41799 25667 41804
rect 23303 41751 23513 41756
rect 5267 40748 5589 40753
rect 218 40436 224 40748
rect 536 40436 5272 40748
rect 5584 40436 5589 40748
rect 5267 40431 5589 40436
rect 5340 37729 5653 37734
rect 3565 37426 3571 37729
rect 3874 37426 5345 37729
rect 5648 37426 5653 37729
rect 5340 37421 5653 37426
<< via3 >>
rect 23306 43916 23506 44116
rect 18252 43308 18452 43508
rect 27038 42990 27238 43190
rect 27580 41804 27780 42004
rect 224 40436 536 40748
rect 3571 37426 3874 37729
<< metal4 >>
rect 200 40748 600 44152
rect 200 40436 224 40748
rect 536 40436 600 40748
rect 200 5740 600 40436
rect 198 5618 600 5740
rect 200 5038 600 5618
rect 198 4966 600 5038
rect 200 1000 600 4966
rect 800 42850 1200 44152
rect 6134 42850 6194 45152
rect 6686 42850 6746 45152
rect 7238 42850 7298 45152
rect 7790 42850 7850 45152
rect 8342 42850 8402 45152
rect 8894 42850 8954 45152
rect 9446 42850 9506 45152
rect 9998 42850 10058 45152
rect 10550 42850 10610 45152
rect 11102 42850 11162 45152
rect 11654 42850 11714 45152
rect 12206 42850 12266 45152
rect 12758 42850 12818 45152
rect 13310 42850 13370 45152
rect 13862 42850 13922 45152
rect 14414 42850 14474 45152
rect 14966 42850 15026 45152
rect 15518 42850 15578 45152
rect 16070 42850 16130 45152
rect 16622 42850 16682 45152
rect 17174 42850 17234 45152
rect 17726 42850 17786 45152
rect 18278 44381 18338 45152
rect 18253 43509 18451 44381
rect 18830 44368 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 18818 44086 18958 44368
rect 23305 44116 23507 44117
rect 23305 44086 23306 44116
rect 18818 43946 23306 44086
rect 23305 43916 23306 43946
rect 23506 43916 23507 44116
rect 27110 43916 27170 45152
rect 23305 43915 23507 43916
rect 18251 43508 18453 43509
rect 18251 43308 18252 43508
rect 18452 43308 18453 43508
rect 18251 43307 18453 43308
rect 27038 43191 27238 43916
rect 27662 43914 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27037 43190 27239 43191
rect 27037 42990 27038 43190
rect 27238 42990 27239 43190
rect 27037 42989 27239 42990
rect 800 42450 17826 42850
rect 800 37729 1200 42450
rect 27598 42005 27763 43914
rect 27579 42004 27781 42005
rect 27579 41804 27580 42004
rect 27780 41804 27781 42004
rect 27579 41803 27781 41804
rect 3570 37729 3875 37730
rect 800 37426 3571 37729
rect 3874 37426 3875 37729
rect 800 1000 1200 37426
rect 3570 37425 3875 37426
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 192
rect 14906 0 15086 192
rect 18770 0 18950 204
rect 22634 0 22814 192
rect 26498 0 26678 200
rect 30362 0 30542 196
use sr_latch  sr_latch_0
timestamp 1770730625
transform 1 0 18026 0 1 42425
box 862 -5005 12821 -1677
use zedulo_logo  zedulo_logo_0 ~/tt_09analog_course/art
timestamp 1771425041
transform 1 0 11638 0 1 15774
box 720 990 8190 7920
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
