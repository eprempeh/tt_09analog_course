magic
tech sky130A
timestamp 1771425041
<< metal4 >>
rect 2655 3915 2880 3960
rect 2745 3870 3015 3915
rect 2835 3825 3105 3870
rect 2925 3780 3195 3825
rect 1215 3735 1260 3780
rect 1620 3735 1755 3780
rect 2970 3735 3285 3780
rect 1035 3690 1350 3735
rect 1395 3690 1485 3735
rect 1710 3690 2025 3735
rect 3015 3690 3420 3735
rect 943 3645 1125 3690
rect 1215 3645 1260 3690
rect 1395 3645 1440 3690
rect 1665 3645 2070 3690
rect 900 3600 990 3645
rect 1350 3600 1440 3645
rect 1620 3600 2070 3645
rect 3060 3645 3465 3690
rect 3060 3600 3510 3645
rect 855 3555 945 3600
rect 1215 3555 1440 3600
rect 1575 3555 2025 3600
rect 3015 3555 3555 3600
rect 810 3510 900 3555
rect 1215 3510 1305 3555
rect 1530 3510 1980 3555
rect 2745 3510 2835 3555
rect 3015 3510 3600 3555
rect 765 3420 855 3510
rect 1035 3420 1125 3510
rect 1440 3465 1935 3510
rect 2745 3465 2790 3510
rect 3015 3465 3645 3510
rect 1395 3420 1845 3465
rect 2970 3420 3690 3465
rect 720 3375 810 3420
rect 900 3375 1125 3420
rect 1350 3375 1620 3420
rect 2970 3375 3735 3420
rect 675 3330 765 3375
rect 855 3330 1080 3375
rect 675 3285 1080 3330
rect 1350 3330 1485 3375
rect 2925 3330 3735 3375
rect 1350 3285 1440 3330
rect 2430 3285 2475 3330
rect 2835 3285 3735 3330
rect 630 3240 1035 3285
rect 1755 3240 1845 3285
rect 585 3195 1035 3240
rect 1800 3195 1845 3240
rect 2340 3240 2655 3285
rect 2790 3240 3780 3285
rect 2340 3195 2700 3240
rect 585 3150 990 3195
rect 540 3060 990 3150
rect 2295 3150 2610 3195
rect 2745 3150 3825 3240
rect 2295 3105 2385 3150
rect 2475 3105 3870 3150
rect 2250 3060 2340 3105
rect 2475 3060 3915 3105
rect 495 2970 810 3060
rect 450 2925 810 2970
rect 450 2880 675 2925
rect 900 2919 952 2971
rect 2205 2925 2340 3060
rect 2430 3015 3915 3060
rect 2475 2970 3960 3015
rect 2520 2925 3960 2970
rect 2250 2880 2295 2925
rect 450 2835 630 2880
rect 450 2790 585 2835
rect 2475 2790 4005 2925
rect 450 2745 540 2790
rect 1935 2745 1980 2790
rect 2430 2745 4050 2790
rect 450 2700 495 2745
rect 1935 2700 2025 2745
rect 2160 2700 4050 2745
rect 2070 2655 4050 2700
rect 2025 2610 4050 2655
rect 1935 2565 3105 2610
rect 1935 2520 3060 2565
rect 3240 2520 4095 2610
rect 360 2340 405 2520
rect 1935 2475 2655 2520
rect 2700 2475 2745 2520
rect 1935 2430 2115 2475
rect 2160 2430 2250 2475
rect 2295 2430 2610 2475
rect 2835 2430 3060 2520
rect 3195 2475 4095 2520
rect 3240 2430 4050 2475
rect 1755 2385 2025 2430
rect 2205 2385 2250 2430
rect 2340 2385 2610 2430
rect 2925 2385 3105 2430
rect 1710 2340 1980 2385
rect 2385 2340 2565 2385
rect 2925 2340 3150 2385
rect 1710 2295 1935 2340
rect 2430 2295 2565 2340
rect 2745 2295 3150 2340
rect 1755 2250 1890 2295
rect 2430 2250 2475 2295
rect 2610 2250 3150 2295
rect 3285 2340 4050 2430
rect 3285 2295 4095 2340
rect 3285 2250 3960 2295
rect 1935 2205 2070 2250
rect 2610 2205 2790 2250
rect 2835 2205 3915 2250
rect 1710 2160 2160 2205
rect 1665 2070 2160 2160
rect 2880 2115 3915 2205
rect 4050 2160 4095 2295
rect 2835 2070 3870 2115
rect 1575 2025 2205 2070
rect 2835 2025 3240 2070
rect 3285 2025 3555 2070
rect 3690 2025 3870 2070
rect 405 1980 450 2025
rect 1530 1980 2250 2025
rect 2430 1980 2520 2025
rect 2700 1980 3240 2025
rect 3735 1980 3870 2025
rect 360 1845 540 1980
rect 1485 1935 3285 1980
rect 1395 1890 2790 1935
rect 2925 1890 3285 1935
rect 3330 1890 3510 1935
rect 3780 1890 3915 1980
rect 4050 1935 4095 1980
rect 360 1800 585 1845
rect 360 1710 630 1800
rect 1395 1755 2835 1890
rect 2925 1845 3465 1890
rect 3015 1755 3465 1845
rect 3825 1800 3870 1890
rect 4005 1845 4095 1935
rect 1395 1710 2880 1755
rect 3060 1710 3420 1755
rect 405 1665 675 1710
rect 1395 1665 2925 1710
rect 405 1575 720 1665
rect 1350 1620 2925 1665
rect 450 1530 720 1575
rect 1395 1575 2925 1620
rect 3105 1665 3375 1710
rect 3105 1620 3330 1665
rect 3105 1575 3240 1620
rect 1395 1530 2970 1575
rect 3150 1530 3195 1575
rect 450 1485 765 1530
rect 1440 1485 3060 1530
rect 495 1395 765 1485
rect 1485 1440 3060 1485
rect 3240 1440 3285 1485
rect 1485 1395 3285 1440
rect 495 1350 810 1395
rect 1575 1350 3285 1395
rect 540 1305 855 1350
rect 585 1260 900 1305
rect 585 1215 990 1260
rect 1431 1257 1488 1310
rect 1665 1305 1755 1350
rect 1845 1305 1890 1350
rect 1935 1305 3240 1350
rect 1980 1260 3195 1305
rect 2115 1215 3150 1260
rect 630 1170 1035 1215
rect 2070 1170 3105 1215
rect 630 1125 1080 1170
rect 2070 1125 3060 1170
rect 3458 1166 3516 1222
rect 675 1080 1125 1125
rect 2115 1080 3015 1125
rect 720 1035 1080 1080
rect 2115 1035 2970 1080
rect 765 945 1080 1035
rect 2205 990 2970 1035
rect 765 900 1035 945
rect 810 855 990 900
rect 1839 894 1905 950
rect 2205 945 2925 990
rect 3015 945 3092 993
rect 3645 945 3690 1035
rect 855 810 990 855
rect 2205 855 2970 945
rect 2205 810 2925 855
rect 900 765 990 810
rect 2160 765 2880 810
rect 3060 765 3150 855
rect 2205 720 2790 765
rect 2250 675 2745 720
rect 1837 581 1914 638
rect 2250 630 2700 675
rect 2250 585 2610 630
rect 2295 540 2565 585
rect 2340 495 2385 540
<< end >>
