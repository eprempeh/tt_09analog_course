magic
tech sky130A
magscale 1 2
timestamp 1771423307
<< metal1 >>
rect 17160 5514 17560 5520
rect 17560 5124 20494 5505
rect 17160 5108 17560 5114
rect 19752 4094 19932 4100
rect 19932 3914 20738 4094
rect 19752 3908 19932 3914
rect 26172 3702 26352 4208
rect 20236 3541 20578 3604
rect 20236 3428 20864 3541
rect 26166 3522 26172 3702
rect 26352 3522 26358 3702
rect 20238 3416 20864 3428
rect 20238 2774 20418 3416
rect 26690 3154 26870 3546
rect 26684 2974 26690 3154
rect 26870 2974 26876 3154
rect 20238 2588 20418 2594
rect 17660 2516 18060 2522
rect 18060 2177 21081 2456
rect 26212 2424 26218 2482
rect 26363 2424 26369 2482
rect 26200 2342 26380 2424
rect 26684 2370 26690 2480
rect 26870 2370 26876 2480
rect 17660 2110 18060 2116
<< via1 >>
rect 17160 5114 17560 5514
rect 19752 3914 19932 4094
rect 26172 3522 26352 3702
rect 26690 2974 26870 3154
rect 20238 2594 20418 2774
rect 17660 2116 18060 2516
<< metal2 >>
rect 14273 5514 14663 5518
rect 14268 5509 17160 5514
rect 14268 5119 14273 5509
rect 14663 5119 17160 5509
rect 14268 5114 17160 5119
rect 17560 5114 17566 5514
rect 14273 5110 14663 5114
rect 19259 4094 19429 4098
rect 19254 4089 19752 4094
rect 19254 3919 19259 4089
rect 19429 3919 19752 4089
rect 19254 3914 19752 3919
rect 19932 3914 19938 4094
rect 19259 3910 19429 3914
rect 26172 3702 26352 3708
rect 26172 3245 26352 3522
rect 26172 3075 26177 3245
rect 26347 3075 26352 3245
rect 26172 3070 26352 3075
rect 26690 3154 26870 3160
rect 26177 3066 26347 3070
rect 26690 2965 26870 2974
rect 26690 2795 26695 2965
rect 26865 2795 26870 2965
rect 26690 2790 26870 2795
rect 26695 2786 26865 2790
rect 20232 2594 20238 2774
rect 20418 2594 20424 2774
rect 16475 2516 16865 2520
rect 16470 2511 17660 2516
rect 16470 2121 16475 2511
rect 16865 2121 17660 2511
rect 16470 2116 17660 2121
rect 18060 2116 18066 2516
rect 16475 2112 16865 2116
rect 20238 1357 20418 2594
rect 20234 1187 20243 1357
rect 20413 1187 20422 1357
rect 20238 1182 20418 1187
<< via2 >>
rect 14273 5119 14663 5509
rect 19259 3919 19429 4089
rect 26177 3075 26347 3245
rect 26695 2795 26865 2965
rect 16475 2121 16865 2511
rect 20243 1187 20413 1357
<< metal3 >>
rect 201 5514 599 5519
rect 200 5513 14668 5514
rect 200 5115 201 5513
rect 599 5509 14668 5513
rect 599 5119 14273 5509
rect 14663 5119 14668 5509
rect 599 5115 14668 5119
rect 200 5114 14668 5115
rect 201 5109 599 5114
rect 18771 4094 18949 4099
rect 18770 4093 19434 4094
rect 18770 3915 18771 4093
rect 18949 4089 19434 4093
rect 18949 3919 19259 4089
rect 19429 3919 19434 4089
rect 18949 3915 19434 3919
rect 18770 3914 19434 3915
rect 18771 3909 18949 3914
rect 26172 3245 26352 3250
rect 26172 3075 26177 3245
rect 26347 3075 26352 3245
rect 12161 2516 12559 2521
rect 12160 2515 16870 2516
rect 12160 2117 12161 2515
rect 12559 2511 16870 2515
rect 12559 2121 16475 2511
rect 16865 2121 16870 2511
rect 12559 2117 16870 2121
rect 12160 2116 16870 2117
rect 12161 2111 12559 2116
rect 26172 1555 26352 3075
rect 26690 2965 26870 2970
rect 26690 2795 26695 2965
rect 26865 2795 26870 2965
rect 26690 1575 26870 2795
rect 26167 1377 26173 1555
rect 26351 1377 26357 1555
rect 26685 1397 26691 1575
rect 26869 1397 26875 1575
rect 26690 1396 26870 1397
rect 26172 1376 26352 1377
rect 20238 1357 20418 1362
rect 20238 1187 20243 1357
rect 20413 1187 20418 1357
rect 20238 755 20418 1187
rect 20233 577 20239 755
rect 20417 577 20423 755
rect 20238 576 20418 577
<< via3 >>
rect 201 5115 599 5513
rect 18771 3915 18949 4093
rect 12161 2117 12559 2515
rect 26173 1377 26351 1555
rect 26691 1397 26869 1575
rect 20239 577 20417 755
<< metal4 >>
rect 200 5513 600 44152
rect 200 5115 201 5513
rect 599 5115 600 5513
rect 200 1000 600 5115
rect 800 42850 1200 44152
rect 6134 42850 6194 45152
rect 6686 42850 6746 45152
rect 7238 42850 7298 45152
rect 7790 42850 7850 45152
rect 8342 42850 8402 45152
rect 8894 42850 8954 45152
rect 9446 42850 9506 45152
rect 9998 42850 10058 45152
rect 10550 42850 10610 45152
rect 11102 42850 11162 45152
rect 11654 42850 11714 45152
rect 12206 42850 12266 45152
rect 12758 42850 12818 45152
rect 13310 42850 13370 45152
rect 13862 42850 13922 45152
rect 14414 42850 14474 45152
rect 14966 42850 15026 45152
rect 15518 42850 15578 45152
rect 16070 42850 16130 45152
rect 16622 42850 16682 45152
rect 17174 42850 17234 45152
rect 17726 42850 17786 45152
rect 18278 42850 18338 45152
rect 18830 42850 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 800 42450 19050 42850
rect 800 2516 1200 42450
rect 18770 4093 18950 4094
rect 18770 3915 18771 4093
rect 18949 3915 18950 4093
rect 800 2515 12560 2516
rect 800 2117 12161 2515
rect 12559 2117 12560 2515
rect 800 2116 12560 2117
rect 800 1000 1200 2116
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 3915
rect 26690 1575 30542 1576
rect 26172 1555 26352 1556
rect 26172 1377 26173 1555
rect 26351 1377 26352 1555
rect 26690 1397 26691 1575
rect 26869 1397 30542 1575
rect 26690 1396 30542 1397
rect 26172 840 26352 1377
rect 20238 755 22814 756
rect 20238 577 20239 755
rect 20417 577 22814 755
rect 26172 660 26678 840
rect 20238 576 22814 577
rect 22634 0 22814 576
rect 26498 0 26678 660
rect 30362 0 30542 1396
use sr_latch  sr_latch_0
timestamp 1770730625
transform 1 0 19230 0 1 7181
box 862 -5005 12821 -1677
use zedulo_logo  zedulo_logo_0 ~/tt_09analog_course/art
timestamp 1771423184
transform 1 0 11774 0 1 19566
box 630 720 8280 8010
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
