magic
tech sky130A
timestamp 1771349514
<< error_p >>
rect 6538 9940 6594 9954
rect 6622 9940 6650 9954
rect 6552 9926 6580 9940
rect 6636 9926 6650 9940
rect 4802 9828 4830 9842
rect 7126 9828 7154 9842
rect 4802 9814 4816 9828
rect 7126 9814 7140 9828
rect 4242 9800 4270 9814
rect 4802 9800 4830 9814
rect 4242 9786 4256 9800
rect 4816 9786 4830 9800
rect 4354 9772 4382 9786
rect 4368 9758 4382 9772
rect 4354 9744 4382 9758
rect 4354 9730 4368 9744
rect 3374 9688 3402 9702
rect 4046 9688 4074 9702
rect 3374 9674 3388 9688
rect 4060 9674 4074 9688
rect 3654 9660 3682 9674
rect 3668 9646 3682 9660
rect 3346 9548 3374 9562
rect 7154 9548 7182 9562
rect 3346 9534 3360 9548
rect 7168 9534 7182 9548
rect 3010 9492 3038 9506
rect 7238 9492 7266 9506
rect 3010 9478 3024 9492
rect 7252 9478 7266 9492
rect 7266 9464 7294 9478
rect 7280 9450 7294 9464
rect 2870 9408 2898 9422
rect 2870 9394 2884 9408
rect 2842 9380 2870 9394
rect 3038 9380 3066 9394
rect 2842 9366 2856 9380
rect 3038 9366 3052 9380
rect 3374 9296 3402 9310
rect 3374 9282 3388 9296
rect 4998 9212 5026 9226
rect 4998 9198 5012 9212
rect 3122 9184 3150 9198
rect 3122 9170 3136 9184
rect 2534 9128 2562 9142
rect 2548 9114 2562 9128
rect 3150 9128 3178 9142
rect 3458 9128 3486 9142
rect 3150 9114 3164 9128
rect 3458 9114 3472 9128
rect 3178 9100 3206 9114
rect 3178 9086 3192 9100
rect 2450 9044 2478 9058
rect 2450 9030 2464 9044
rect 3458 8932 3486 8946
rect 6622 8932 6650 8946
rect 3458 8918 3472 8932
rect 6622 8918 6636 8932
rect 4998 8876 5026 8890
rect 4998 8862 5012 8876
rect 3822 8848 3850 8862
rect 7098 8848 7126 8862
rect 7490 8848 7518 8862
rect 3822 8834 3836 8848
rect 7098 8834 7112 8848
rect 7504 8834 7518 8848
rect 4522 8708 4550 8722
rect 5754 8708 5782 8722
rect 4536 8694 4550 8708
rect 5768 8694 5782 8708
rect 7630 8680 7658 8694
rect 7630 8666 7644 8680
rect 7658 8624 7686 8638
rect 7672 8610 7686 8624
rect 4690 8596 4746 8610
rect 4704 8582 4732 8596
rect 2842 8568 2870 8582
rect 2842 8554 2856 8568
rect 4326 8512 4354 8526
rect 4340 8498 4354 8512
rect 8414 8428 8442 8442
rect 8428 8414 8442 8428
rect 2310 8400 2338 8414
rect 2310 8386 2324 8400
rect 7266 8288 7294 8302
rect 7266 8274 7280 8288
rect 8022 8204 8050 8218
rect 8036 8190 8050 8204
rect 6958 8148 6986 8162
rect 6972 8134 6986 8148
rect 6846 8092 6874 8106
rect 6860 8078 6874 8092
rect 6930 8064 6958 8078
rect 6930 8050 6944 8064
rect 8330 7896 8358 7910
rect 8554 7896 8582 7910
rect 8344 7882 8358 7896
rect 8568 7882 8582 7896
rect 7518 7644 7546 7658
rect 7518 7630 7532 7644
rect 5474 7308 5502 7322
rect 5474 7294 5488 7308
rect 4830 6888 4858 6902
rect 4830 6874 4844 6888
rect 938 6832 966 6846
rect 938 6818 952 6832
rect 5222 6748 5250 6762
rect 5222 6734 5236 6748
rect 6510 6132 6538 6146
rect 6510 6118 6524 6132
rect 4970 6048 4998 6062
rect 4970 6034 4984 6048
rect 5446 6020 5474 6034
rect 5460 6006 5474 6020
rect 5642 5852 5670 5866
rect 5656 5838 5670 5852
rect 10150 5852 10178 5866
rect 10150 5838 10164 5852
rect 5306 5712 5334 5726
rect 5306 5698 5320 5712
rect 9450 5628 9478 5642
rect 9464 5614 9478 5628
rect 6510 5544 6538 5558
rect 6524 5530 6538 5544
rect 4046 5124 4074 5138
rect 4046 5110 4060 5124
rect 6118 5068 6146 5082
rect 6132 5054 6146 5068
rect 6874 5040 6902 5054
rect 8190 5040 8218 5054
rect 6888 5026 6902 5040
rect 8204 5026 8218 5040
rect 8218 5012 8246 5026
rect 8232 4998 8246 5012
rect 3878 4984 3906 4998
rect 3878 4970 3892 4984
rect 686 4452 714 4466
rect 686 4438 700 4452
rect 1470 4424 1498 4438
rect 1484 4410 1498 4424
rect 1134 4284 1162 4298
rect 1134 4270 1148 4284
rect 8386 4228 8414 4242
rect 8386 4214 8400 4228
rect 1638 4172 1666 4186
rect 1652 4158 1666 4172
rect 3598 3724 3626 3738
rect 3612 3710 3626 3724
rect 3626 3696 3654 3710
rect 3640 3682 3654 3696
rect 7714 3612 7742 3626
rect 7728 3598 7742 3612
rect 5166 2828 5194 2842
rect 5180 2814 5194 2828
rect 2366 2688 2394 2702
rect 2366 2674 2380 2688
rect 2450 2212 2478 2226
rect 2450 2198 2464 2212
<< metal2 >>
rect 5040 10360 5068 10388
rect 7028 10136 7056 10164
rect 5852 10024 5880 10052
rect 5936 10024 5992 10052
rect 6468 9912 6496 9968
rect 6524 9940 6552 9968
rect 6580 9940 6636 9968
rect 6944 9940 6972 9968
rect 6552 9912 6580 9940
rect 6636 9912 6748 9940
rect 6944 9912 7028 9940
rect 6524 9884 6580 9912
rect 6608 9884 6748 9912
rect 6776 9884 6832 9912
rect 7056 9884 7112 9912
rect 6608 9856 6916 9884
rect 7084 9856 7224 9884
rect 8232 9856 8288 9884
rect 3136 9828 3164 9856
rect 4816 9828 4844 9856
rect 4872 9828 4928 9856
rect 6664 9828 7028 9856
rect 7140 9828 7168 9856
rect 7196 9828 7280 9856
rect 8232 9828 8260 9856
rect 3640 9800 3696 9828
rect 4256 9800 4312 9828
rect 4704 9800 4816 9828
rect 4900 9800 5012 9828
rect 6524 9800 6608 9828
rect 6636 9800 7084 9828
rect 7112 9800 7140 9828
rect 7224 9800 7364 9828
rect 3584 9772 3612 9800
rect 4060 9772 4088 9800
rect 3500 9744 3528 9772
rect 4032 9744 4144 9772
rect 4228 9744 4256 9800
rect 4284 9772 4368 9800
rect 4816 9772 4872 9800
rect 6552 9772 6692 9800
rect 6776 9772 7168 9800
rect 7252 9772 7420 9800
rect 7896 9772 7924 9800
rect 4368 9744 4396 9772
rect 4536 9744 4704 9772
rect 4760 9744 4788 9772
rect 6804 9744 7476 9772
rect 4088 9716 4116 9744
rect 4228 9716 4284 9744
rect 3388 9688 3444 9716
rect 3640 9688 3752 9716
rect 4032 9688 4060 9716
rect 4340 9688 4368 9744
rect 4536 9716 4676 9744
rect 6832 9716 7364 9744
rect 7392 9716 7532 9744
rect 3332 9660 3388 9688
rect 3472 9660 3500 9688
rect 3640 9660 3668 9688
rect 4060 9660 4116 9688
rect 4312 9660 4368 9688
rect 4480 9688 4592 9716
rect 6860 9688 7420 9716
rect 7448 9688 7588 9716
rect 4480 9660 4508 9688
rect 6916 9660 7644 9688
rect 3304 9632 3360 9660
rect 3668 9632 3752 9660
rect 3808 9632 3836 9660
rect 4060 9632 4088 9660
rect 6944 9632 7728 9660
rect 3220 9604 3276 9632
rect 3668 9604 3696 9632
rect 3780 9604 3864 9632
rect 4368 9604 4452 9632
rect 6972 9604 7756 9632
rect 3192 9576 3248 9604
rect 3668 9576 3836 9604
rect 4284 9576 4424 9604
rect 7084 9576 7168 9604
rect 7196 9576 7812 9604
rect 3108 9548 3164 9576
rect 3360 9548 3416 9576
rect 3584 9548 3640 9576
rect 3724 9548 3780 9576
rect 3892 9548 3948 9576
rect 4172 9548 4228 9576
rect 4312 9548 4396 9576
rect 4452 9548 4508 9576
rect 7112 9548 7168 9576
rect 7280 9548 7868 9576
rect 3052 9520 3136 9548
rect 3304 9520 3360 9548
rect 3388 9520 3444 9548
rect 3472 9520 3640 9548
rect 3864 9520 4004 9548
rect 4144 9520 4256 9548
rect 4368 9520 4508 9548
rect 7168 9520 7224 9548
rect 7336 9520 7924 9548
rect 2660 9492 2688 9520
rect 3024 9492 3080 9520
rect 3108 9492 3136 9520
rect 3416 9492 3444 9520
rect 3528 9492 3612 9520
rect 3864 9492 3948 9520
rect 4060 9492 4116 9520
rect 4424 9492 4452 9520
rect 7196 9492 7252 9520
rect 7364 9492 7952 9520
rect 2968 9464 3024 9492
rect 3780 9464 3836 9492
rect 4032 9464 4116 9492
rect 4284 9464 4312 9492
rect 7252 9464 7280 9492
rect 7392 9464 8008 9492
rect 3052 9436 3080 9464
rect 3948 9436 4060 9464
rect 4088 9436 4144 9464
rect 4200 9436 4368 9464
rect 6776 9436 6832 9464
rect 7028 9436 7056 9464
rect 7280 9436 7336 9464
rect 7448 9436 8064 9464
rect 2884 9408 2912 9436
rect 3920 9408 4396 9436
rect 7000 9408 7140 9436
rect 7364 9408 8120 9436
rect 2856 9380 2884 9408
rect 3052 9380 3080 9408
rect 3192 9380 3248 9408
rect 3444 9380 3556 9408
rect 3640 9380 3780 9408
rect 3976 9380 4256 9408
rect 7056 9380 7112 9408
rect 7420 9380 8148 9408
rect 2800 9352 2856 9380
rect 2968 9352 3052 9380
rect 3108 9352 3220 9380
rect 3332 9352 3500 9380
rect 3612 9352 3808 9380
rect 4004 9352 4284 9380
rect 4312 9352 4340 9380
rect 4424 9352 4704 9380
rect 7476 9352 8176 9380
rect 2772 9296 2828 9352
rect 2940 9324 3024 9352
rect 3080 9324 3192 9352
rect 3304 9324 3444 9352
rect 3556 9324 3808 9352
rect 4228 9324 4816 9352
rect 7448 9324 8232 9352
rect 2912 9296 2996 9324
rect 3080 9296 3164 9324
rect 3304 9296 3360 9324
rect 3388 9296 3416 9324
rect 3500 9296 3780 9324
rect 4228 9296 4396 9324
rect 4424 9296 4536 9324
rect 4564 9296 4620 9324
rect 4648 9296 4676 9324
rect 4732 9296 4956 9324
rect 7476 9296 8288 9324
rect 2688 9268 2716 9296
rect 2912 9268 2968 9296
rect 3052 9268 3136 9296
rect 3276 9268 3388 9296
rect 3472 9268 3780 9296
rect 4256 9268 4760 9296
rect 4788 9268 4984 9296
rect 7504 9268 8316 9296
rect 2632 9240 2660 9268
rect 2744 9240 2772 9268
rect 2884 9240 2996 9268
rect 3024 9240 3108 9268
rect 3220 9240 3388 9268
rect 3444 9240 3780 9268
rect 4200 9240 4312 9268
rect 4340 9240 5040 9268
rect 7224 9240 7364 9268
rect 7532 9240 8344 9268
rect 8708 9240 8736 9268
rect 2604 9212 2660 9240
rect 2800 9212 3052 9240
rect 3164 9212 3360 9240
rect 3444 9212 3752 9240
rect 2548 9184 2632 9212
rect 2520 9156 2604 9184
rect 2716 9156 2744 9212
rect 2800 9184 2856 9212
rect 2884 9184 2996 9212
rect 3136 9184 3360 9212
rect 3472 9184 3752 9212
rect 4228 9212 4984 9240
rect 5012 9212 5040 9240
rect 7280 9212 7448 9240
rect 7588 9212 8400 9240
rect 8680 9212 8736 9240
rect 4228 9184 4368 9212
rect 4396 9184 4732 9212
rect 4760 9184 5012 9212
rect 7364 9184 7560 9212
rect 7644 9184 8428 9212
rect 2772 9156 2912 9184
rect 3080 9156 3136 9184
rect 2492 9128 2548 9156
rect 2688 9128 2856 9156
rect 3052 9128 3136 9156
rect 3164 9156 3332 9184
rect 3164 9128 3304 9156
rect 3472 9128 3696 9184
rect 4200 9156 4452 9184
rect 4480 9156 5040 9184
rect 7504 9156 8456 9184
rect 4200 9128 5152 9156
rect 7504 9128 8512 9156
rect 2464 9100 2520 9128
rect 2408 9072 2520 9100
rect 2548 9072 2632 9128
rect 2688 9100 2744 9128
rect 2996 9100 3164 9128
rect 3192 9100 3304 9128
rect 3444 9100 3472 9128
rect 3500 9100 3640 9128
rect 4172 9100 4340 9128
rect 4368 9100 4648 9128
rect 4676 9100 4928 9128
rect 4956 9100 5068 9128
rect 7560 9100 8540 9128
rect 2660 9072 2744 9100
rect 2856 9072 2912 9100
rect 2968 9072 3192 9100
rect 3444 9072 3612 9100
rect 4144 9072 4424 9100
rect 4452 9072 4704 9100
rect 4732 9072 5068 9100
rect 2072 9044 2100 9072
rect 2380 9044 2436 9072
rect 2464 9044 2492 9072
rect 2352 9016 2464 9044
rect 2548 9016 2604 9072
rect 2660 9016 2716 9072
rect 2772 9044 2912 9072
rect 3052 9044 3164 9072
rect 3416 9044 3584 9072
rect 4116 9044 4480 9072
rect 4508 9044 4788 9072
rect 4816 9044 5152 9072
rect 7224 9044 7252 9100
rect 7560 9072 8568 9100
rect 7560 9044 8596 9072
rect 2744 9016 2912 9044
rect 3024 9016 3108 9044
rect 3388 9016 3556 9044
rect 3948 9016 4032 9044
rect 4060 9016 4256 9044
rect 4284 9016 4564 9044
rect 4592 9016 4956 9044
rect 4984 9016 5180 9044
rect 7560 9016 7616 9044
rect 7644 9016 8652 9044
rect 8848 9016 8904 9044
rect 2324 8988 2492 9016
rect 2296 8960 2408 8988
rect 1988 8932 2044 8960
rect 2268 8932 2380 8960
rect 1988 8904 2072 8932
rect 2240 8904 2324 8932
rect 2044 8876 2072 8904
rect 2184 8876 2296 8904
rect 2156 8848 2296 8876
rect 2128 8820 2296 8848
rect 2100 8792 2240 8820
rect 2072 8764 2212 8792
rect 2268 8764 2296 8820
rect 2352 8792 2380 8932
rect 2436 8904 2464 8988
rect 2520 8932 2576 9016
rect 2632 8988 2688 9016
rect 2744 8988 2884 9016
rect 2968 8988 3052 9016
rect 3332 8988 3500 9016
rect 3976 8988 4144 9016
rect 4172 8988 5068 9016
rect 5124 8988 5264 9016
rect 6552 8988 6692 9016
rect 2940 8960 2996 8988
rect 3304 8960 3500 8988
rect 4004 8960 4424 8988
rect 4480 8960 4648 8988
rect 4676 8960 5152 8988
rect 6496 8960 6692 8988
rect 7588 8988 8680 9016
rect 7588 8960 8708 8988
rect 3332 8932 3444 8960
rect 3472 8932 3528 8960
rect 4004 8932 4200 8960
rect 4228 8932 4508 8960
rect 4564 8932 4816 8960
rect 4844 8932 5152 8960
rect 6440 8932 6468 8960
rect 6496 8932 6552 8960
rect 6636 8932 6692 8960
rect 7644 8932 8736 8960
rect 2520 8876 2548 8932
rect 3276 8904 3472 8932
rect 3976 8904 4928 8932
rect 3052 8876 3080 8904
rect 3108 8876 3472 8904
rect 3948 8876 4060 8904
rect 4088 8876 4396 8904
rect 2828 8848 2856 8876
rect 3024 8848 3472 8876
rect 3836 8848 3864 8876
rect 3948 8848 4172 8876
rect 4200 8848 4396 8876
rect 4424 8848 4704 8904
rect 4732 8876 4928 8904
rect 5012 8876 5040 8932
rect 6440 8904 6636 8932
rect 7084 8904 7112 8932
rect 7532 8904 8764 8932
rect 6440 8876 6580 8904
rect 7056 8876 7140 8904
rect 4732 8848 4788 8876
rect 2772 8820 2856 8848
rect 2968 8820 3332 8848
rect 3360 8820 3472 8848
rect 3808 8820 3836 8848
rect 3920 8820 4480 8848
rect 4508 8820 4564 8848
rect 2940 8792 3304 8820
rect 3360 8792 3444 8820
rect 3892 8792 3948 8820
rect 4004 8792 4284 8820
rect 4312 8792 4564 8820
rect 4592 8820 4788 8848
rect 4816 8848 5012 8876
rect 7000 8848 7084 8876
rect 7112 8848 7140 8876
rect 7476 8848 7504 8904
rect 7532 8876 8792 8904
rect 7532 8848 8820 8876
rect 4816 8820 4872 8848
rect 4928 8820 4956 8848
rect 5796 8820 5824 8848
rect 5936 8820 5964 8848
rect 6972 8820 7112 8848
rect 7504 8820 8848 8848
rect 4592 8792 4648 8820
rect 2940 8764 3192 8792
rect 3220 8764 3276 8792
rect 3864 8764 4032 8792
rect 4060 8764 4340 8792
rect 4368 8764 4648 8792
rect 4676 8792 4872 8820
rect 5684 8792 5740 8820
rect 5796 8792 5852 8820
rect 5880 8792 5992 8820
rect 6916 8792 7084 8820
rect 7532 8792 8876 8820
rect 4676 8764 4900 8792
rect 5712 8764 5992 8792
rect 6888 8764 7028 8792
rect 7532 8764 8904 8792
rect 2044 8736 2212 8764
rect 2240 8736 2296 8764
rect 1680 8708 1736 8736
rect 2016 8708 2212 8736
rect 1988 8652 2128 8708
rect 1708 8624 1736 8652
rect 1932 8624 2128 8652
rect 1904 8568 2128 8624
rect 1596 8540 1624 8568
rect 1876 8540 2128 8568
rect 1708 8484 1736 8540
rect 1848 8512 2044 8540
rect 1820 8456 2044 8512
rect 1540 8428 1568 8456
rect 1792 8428 1960 8456
rect 1764 8400 1960 8428
rect 1736 8372 1960 8400
rect 1708 8316 1960 8372
rect 1680 8288 1960 8316
rect 1988 8288 2044 8456
rect 2072 8484 2128 8540
rect 2156 8540 2212 8708
rect 2324 8680 2352 8764
rect 3052 8736 3136 8764
rect 3220 8736 3248 8764
rect 3724 8736 3808 8764
rect 2716 8680 2800 8708
rect 3024 8680 3136 8736
rect 3192 8708 3248 8736
rect 3696 8708 3808 8736
rect 3836 8736 4424 8764
rect 4480 8736 4732 8764
rect 4760 8736 4956 8764
rect 5740 8736 5880 8764
rect 6860 8736 7028 8764
rect 7560 8736 7616 8764
rect 7644 8736 8932 8764
rect 3836 8708 4116 8736
rect 4172 8708 4536 8736
rect 4564 8708 4844 8736
rect 5740 8708 5768 8736
rect 5824 8708 5908 8736
rect 3220 8680 3248 8708
rect 3584 8680 3920 8708
rect 3948 8680 4200 8708
rect 4228 8680 4508 8708
rect 4536 8680 4592 8708
rect 4648 8680 4844 8708
rect 5768 8680 5880 8708
rect 6888 8680 7000 8736
rect 7560 8708 8960 8736
rect 7504 8680 7616 8708
rect 7644 8680 7700 8708
rect 7756 8680 8988 8708
rect 2240 8596 2268 8680
rect 2688 8652 2828 8680
rect 2632 8624 2828 8652
rect 2996 8624 3136 8680
rect 3584 8652 3724 8680
rect 3752 8652 4284 8680
rect 4312 8652 4704 8680
rect 3556 8624 4368 8652
rect 4424 8624 4676 8652
rect 4732 8624 4788 8680
rect 5796 8652 5880 8680
rect 5824 8624 5880 8652
rect 6860 8652 7000 8680
rect 7252 8652 7308 8680
rect 7420 8652 7644 8680
rect 7784 8652 9016 8680
rect 6860 8624 6888 8652
rect 2604 8568 2828 8624
rect 2856 8568 2884 8624
rect 2996 8596 3080 8624
rect 3528 8596 3836 8624
rect 3024 8568 3052 8596
rect 3472 8568 3584 8596
rect 3612 8568 3836 8596
rect 3864 8596 4452 8624
rect 4508 8596 4704 8624
rect 4732 8596 4760 8624
rect 6860 8596 6916 8624
rect 6944 8596 7000 8652
rect 3864 8568 4144 8596
rect 4200 8568 4536 8596
rect 4592 8568 4648 8596
rect 4704 8568 4732 8596
rect 2576 8540 2856 8568
rect 2156 8512 2184 8540
rect 2520 8512 2856 8540
rect 3472 8540 3640 8568
rect 3668 8540 4228 8568
rect 4284 8540 4620 8568
rect 6860 8540 7000 8596
rect 7280 8624 7364 8652
rect 7420 8624 7672 8652
rect 7784 8624 9044 8652
rect 9268 8624 9296 8652
rect 7280 8596 7392 8624
rect 7448 8596 7644 8624
rect 7672 8596 7700 8624
rect 7756 8596 8484 8624
rect 8512 8596 9072 8624
rect 7280 8568 7420 8596
rect 7476 8568 7532 8596
rect 7560 8568 7644 8596
rect 7728 8568 9100 8596
rect 7308 8540 7448 8568
rect 7560 8540 7672 8568
rect 7700 8540 8036 8568
rect 8064 8540 9128 8568
rect 3472 8512 3920 8540
rect 3948 8512 4340 8540
rect 4368 8512 4648 8540
rect 6860 8512 6944 8540
rect 2408 8484 2436 8512
rect 2464 8484 2492 8512
rect 2520 8484 2716 8512
rect 2744 8484 2884 8512
rect 3444 8484 3500 8512
rect 3528 8484 4032 8512
rect 4060 8484 4312 8512
rect 4340 8484 4396 8512
rect 4592 8484 4620 8512
rect 5152 8484 5180 8512
rect 6888 8484 6944 8512
rect 6972 8512 7000 8540
rect 7336 8512 7476 8540
rect 7560 8512 7812 8540
rect 7840 8512 9156 8540
rect 6972 8484 7028 8512
rect 2072 8428 2100 8484
rect 2268 8456 2296 8484
rect 2352 8456 2884 8484
rect 2324 8428 2884 8456
rect 3416 8456 3780 8484
rect 3808 8456 4116 8484
rect 4144 8456 4368 8484
rect 6888 8456 7056 8484
rect 7392 8456 7532 8512
rect 7560 8484 8288 8512
rect 8316 8484 8456 8512
rect 8484 8484 8596 8512
rect 8624 8484 9184 8512
rect 9464 8484 9492 8512
rect 7588 8456 7728 8484
rect 7784 8456 7952 8484
rect 7980 8456 8120 8484
rect 8148 8456 9184 8484
rect 3416 8428 3864 8456
rect 3892 8428 4172 8456
rect 4228 8428 4452 8456
rect 6300 8428 6328 8456
rect 7000 8428 7112 8456
rect 7168 8428 7280 8456
rect 2072 8400 2128 8428
rect 2100 8288 2128 8400
rect 2184 8372 2212 8428
rect 2324 8400 2548 8428
rect 2576 8400 2716 8428
rect 2744 8400 2800 8428
rect 3388 8400 3948 8428
rect 3976 8400 4004 8428
rect 4312 8400 4564 8428
rect 7196 8400 7364 8428
rect 7448 8400 7560 8456
rect 7616 8428 8260 8456
rect 7700 8400 8064 8428
rect 8092 8400 8260 8428
rect 8288 8428 8428 8456
rect 8456 8428 9212 8456
rect 8288 8400 8400 8428
rect 8428 8400 8568 8428
rect 8596 8400 9240 8428
rect 2268 8372 2324 8400
rect 2352 8372 2688 8400
rect 2744 8372 2772 8400
rect 3360 8372 3444 8400
rect 3472 8372 3948 8400
rect 4424 8372 4480 8400
rect 4508 8372 4564 8400
rect 7504 8372 7588 8400
rect 7644 8372 9268 8400
rect 9464 8372 9520 8400
rect 2240 8344 2660 8372
rect 3360 8344 3808 8372
rect 3836 8344 3948 8372
rect 7392 8344 7448 8372
rect 7476 8344 7616 8372
rect 2212 8316 2688 8344
rect 2716 8316 2744 8344
rect 3332 8316 3556 8344
rect 3584 8316 3780 8344
rect 7308 8316 7364 8344
rect 2156 8288 2688 8316
rect 2912 8288 2940 8316
rect 3332 8288 3360 8316
rect 3388 8288 3696 8316
rect 7196 8288 7252 8316
rect 7280 8288 7364 8316
rect 1652 8260 1960 8288
rect 2016 8260 2044 8288
rect 2156 8260 2716 8288
rect 3332 8260 3640 8288
rect 7112 8260 7280 8288
rect 1624 8232 1960 8260
rect 1596 8176 1960 8232
rect 2128 8232 2716 8260
rect 3304 8232 3444 8260
rect 3472 8232 3612 8260
rect 6076 8232 6216 8260
rect 7056 8232 7196 8260
rect 2128 8204 2688 8232
rect 3304 8204 3584 8232
rect 6076 8204 6300 8232
rect 7028 8204 7196 8232
rect 7224 8232 7280 8260
rect 7308 8260 7364 8288
rect 7392 8316 7532 8344
rect 7588 8316 7616 8344
rect 7672 8344 7812 8372
rect 7840 8344 8008 8372
rect 8036 8344 8204 8372
rect 8232 8344 9296 8372
rect 9464 8344 9492 8372
rect 7672 8316 7728 8344
rect 7784 8316 7952 8344
rect 7980 8316 8148 8344
rect 7392 8288 7644 8316
rect 7392 8260 7588 8288
rect 7308 8232 7588 8260
rect 7616 8260 7644 8288
rect 7700 8288 8148 8316
rect 8176 8316 8344 8344
rect 8400 8316 8512 8344
rect 8176 8288 8512 8316
rect 8540 8316 9296 8344
rect 8540 8288 9324 8316
rect 7700 8260 7896 8288
rect 7924 8260 8092 8288
rect 8120 8260 8316 8288
rect 8344 8260 8792 8288
rect 8820 8260 9352 8288
rect 7616 8232 7812 8260
rect 7224 8204 7448 8232
rect 7476 8204 7532 8232
rect 7560 8204 7812 8232
rect 7840 8232 8232 8260
rect 7840 8204 8036 8232
rect 8064 8204 8232 8232
rect 8288 8232 8456 8260
rect 8512 8232 8624 8260
rect 8288 8204 8624 8232
rect 8652 8232 9380 8260
rect 8652 8204 9408 8232
rect 2072 8176 2660 8204
rect 3276 8176 3528 8204
rect 1568 8148 1988 8176
rect 2044 8148 2660 8176
rect 3304 8148 3332 8176
rect 3360 8148 3500 8176
rect 4088 8148 4116 8176
rect 4368 8148 4424 8204
rect 5936 8176 5964 8204
rect 6048 8176 6328 8204
rect 5908 8148 6328 8176
rect 6384 8148 6440 8176
rect 1540 8120 1904 8148
rect 1932 8120 2016 8148
rect 1512 8092 2016 8120
rect 2044 8092 2632 8148
rect 3360 8120 3444 8148
rect 4368 8120 4452 8148
rect 5880 8120 6048 8148
rect 3388 8092 3416 8120
rect 4340 8092 4452 8120
rect 4480 8092 4564 8120
rect 4592 8092 4648 8120
rect 1512 8064 2632 8092
rect 1484 8036 2632 8064
rect 4368 8036 4648 8092
rect 5880 8092 5936 8120
rect 5992 8092 6048 8120
rect 6076 8120 6216 8148
rect 6272 8120 6440 8148
rect 6076 8092 6132 8120
rect 5880 8064 6132 8092
rect 6188 8092 6244 8120
rect 6272 8092 6328 8120
rect 6356 8092 6440 8120
rect 6468 8148 6524 8176
rect 6468 8092 6552 8148
rect 6804 8120 6860 8176
rect 6944 8148 6972 8204
rect 7028 8176 7084 8204
rect 7112 8176 7420 8204
rect 7476 8176 7728 8204
rect 7784 8176 8008 8204
rect 8036 8176 8400 8204
rect 8456 8176 9408 8204
rect 9744 8176 9772 8204
rect 7028 8148 7336 8176
rect 7364 8148 7672 8176
rect 7700 8148 7952 8176
rect 7980 8148 8176 8176
rect 8204 8148 8568 8176
rect 8624 8148 8736 8176
rect 8764 8148 9436 8176
rect 6580 8092 6664 8120
rect 6832 8092 6860 8120
rect 6972 8120 7000 8148
rect 7028 8120 7252 8148
rect 6972 8092 7140 8120
rect 6188 8064 6692 8092
rect 5824 8036 6580 8064
rect 1456 8008 2604 8036
rect 4340 8008 4480 8036
rect 1456 7980 2436 8008
rect 1428 7952 2436 7980
rect 2464 7980 2576 8008
rect 4368 7980 4480 8008
rect 4508 8008 4676 8036
rect 5824 8008 6272 8036
rect 4508 7980 4648 8008
rect 5488 7980 5544 8008
rect 2464 7952 2548 7980
rect 4368 7952 4564 7980
rect 5824 7952 5880 8008
rect 5908 7980 5964 8008
rect 5992 7980 6048 8008
rect 6104 7980 6160 8008
rect 6216 7980 6272 8008
rect 6300 7980 6384 8036
rect 6412 8008 6468 8036
rect 6524 8008 6580 8036
rect 6636 8036 6692 8064
rect 6720 8036 6776 8064
rect 6860 8036 6888 8092
rect 6944 8064 7056 8092
rect 6636 8008 6776 8036
rect 6916 8008 6944 8064
rect 7000 8036 7056 8064
rect 7084 8064 7140 8092
rect 7168 8092 7252 8120
rect 7280 8120 7588 8148
rect 7616 8120 7868 8148
rect 7924 8120 8120 8148
rect 7280 8092 7560 8120
rect 7616 8092 7812 8120
rect 7168 8064 7476 8092
rect 7532 8064 7812 8092
rect 7840 8092 8120 8120
rect 8148 8120 8344 8148
rect 8400 8120 8904 8148
rect 8932 8120 9464 8148
rect 8148 8092 9464 8120
rect 7840 8064 8036 8092
rect 8092 8064 8288 8092
rect 7084 8036 7392 8064
rect 7448 8036 7728 8064
rect 7784 8036 7980 8064
rect 8008 8036 8288 8064
rect 8316 8064 8512 8092
rect 8568 8064 8680 8092
rect 8736 8064 8848 8092
rect 8904 8064 9492 8092
rect 8316 8036 8708 8064
rect 8736 8036 8876 8064
rect 8904 8036 9520 8064
rect 7000 8008 7280 8036
rect 7336 8008 7644 8036
rect 6412 7980 6776 8008
rect 6860 7980 7196 8008
rect 5908 7952 6692 7980
rect 6832 7952 7112 7980
rect 7140 7952 7196 7980
rect 7224 7980 7308 8008
rect 7336 7980 7560 8008
rect 7588 7980 7644 8008
rect 7672 8008 7952 8036
rect 8008 8008 8204 8036
rect 8232 8008 8484 8036
rect 8512 8008 9548 8036
rect 9716 8008 9772 8064
rect 7672 7980 7896 8008
rect 7224 7952 7532 7980
rect 7588 7952 7896 7980
rect 7924 7980 8428 8008
rect 7924 7952 8120 7980
rect 8176 7952 8428 7980
rect 8456 7980 8624 8008
rect 8680 7980 8988 8008
rect 9016 7980 9548 8008
rect 9744 7980 9772 8008
rect 8456 7952 8652 7980
rect 8680 7952 8820 7980
rect 8848 7952 9548 7980
rect 1428 7924 2576 7952
rect 4452 7924 4480 7952
rect 5796 7924 6412 7952
rect 1400 7896 2520 7924
rect 2548 7896 2576 7924
rect 5796 7896 5992 7924
rect 1372 7868 2520 7896
rect 5768 7868 5880 7896
rect 5936 7868 5992 7896
rect 6020 7896 6104 7924
rect 6132 7896 6188 7924
rect 6020 7868 6076 7896
rect 6160 7868 6188 7896
rect 6216 7896 6300 7924
rect 6328 7896 6412 7924
rect 6440 7924 6496 7952
rect 6804 7924 7000 7952
rect 7028 7924 7084 7952
rect 7140 7924 7448 7952
rect 6440 7896 6524 7924
rect 6804 7896 6888 7924
rect 6216 7868 6524 7896
rect 6720 7868 6748 7896
rect 1372 7840 2548 7868
rect 1176 7812 1204 7840
rect 1344 7784 2548 7840
rect 5740 7812 6076 7868
rect 3416 7784 3444 7812
rect 1316 7728 2548 7784
rect 4648 7756 4676 7784
rect 5040 7756 5068 7784
rect 5684 7756 5712 7784
rect 5740 7756 5796 7812
rect 5852 7756 5908 7812
rect 5936 7784 6076 7812
rect 6216 7840 6552 7868
rect 6692 7840 6748 7868
rect 6832 7868 6888 7896
rect 6916 7896 6972 7924
rect 7028 7896 7364 7924
rect 6916 7868 7252 7896
rect 7280 7868 7364 7896
rect 7392 7896 7448 7924
rect 7504 7924 7784 7952
rect 7840 7924 8344 7952
rect 7504 7896 7700 7924
rect 7392 7868 7700 7896
rect 7756 7896 8064 7924
rect 8092 7896 8232 7924
rect 8316 7896 8344 7924
rect 8372 7924 8596 7952
rect 8624 7924 9576 7952
rect 8372 7896 8568 7924
rect 8652 7896 8960 7924
rect 8988 7896 9604 7924
rect 7756 7868 7952 7896
rect 6832 7840 7252 7868
rect 7308 7840 7616 7868
rect 7672 7840 7952 7868
rect 8008 7840 8232 7896
rect 8344 7840 8512 7896
rect 8568 7868 8764 7896
rect 8792 7868 9100 7896
rect 9128 7868 9632 7896
rect 8568 7840 9632 7868
rect 6216 7812 6440 7840
rect 6216 7784 6328 7812
rect 6384 7784 6440 7812
rect 6496 7784 6552 7840
rect 6720 7812 7028 7840
rect 6748 7784 7028 7812
rect 7084 7812 7140 7840
rect 7196 7812 7532 7840
rect 7588 7812 7868 7840
rect 7924 7812 8260 7840
rect 8288 7812 8456 7840
rect 8484 7812 8708 7840
rect 8736 7812 8932 7840
rect 8960 7812 9072 7840
rect 7084 7784 7420 7812
rect 5936 7756 6020 7784
rect 6244 7756 6692 7784
rect 6720 7756 6804 7784
rect 6860 7756 6916 7784
rect 6972 7756 7308 7784
rect 1288 7700 2548 7728
rect 3556 7700 3584 7756
rect 3976 7728 4004 7756
rect 5656 7728 6020 7756
rect 6188 7728 6608 7756
rect 6636 7728 6692 7756
rect 6748 7728 6832 7756
rect 6860 7728 7168 7756
rect 5628 7700 6020 7728
rect 6132 7700 6496 7728
rect 6524 7700 6580 7728
rect 6636 7700 7168 7728
rect 7252 7700 7308 7756
rect 7364 7756 7420 7784
rect 7476 7784 7532 7812
rect 7560 7784 7784 7812
rect 7476 7756 7784 7784
rect 7840 7784 7896 7812
rect 7924 7784 8120 7812
rect 7840 7756 8120 7784
rect 8176 7784 8456 7812
rect 8512 7784 9072 7812
rect 9100 7784 9660 7840
rect 8176 7756 8372 7784
rect 7364 7728 7700 7756
rect 7756 7728 8036 7756
rect 8092 7728 8372 7756
rect 8428 7756 8652 7784
rect 8708 7756 8876 7784
rect 8904 7756 9688 7784
rect 8428 7728 9044 7756
rect 9072 7728 9688 7756
rect 7364 7700 7588 7728
rect 1092 7672 1120 7700
rect 1288 7672 2100 7700
rect 2156 7672 2520 7700
rect 5404 7672 5432 7700
rect 1260 7616 1372 7672
rect 1232 7588 1372 7616
rect 1204 7560 1372 7588
rect 1456 7644 2100 7672
rect 2184 7644 2520 7672
rect 3276 7644 3332 7672
rect 1456 7616 2072 7644
rect 2184 7616 2464 7644
rect 3248 7616 3332 7644
rect 5572 7644 5712 7700
rect 5740 7644 5796 7700
rect 5852 7644 5908 7700
rect 6188 7672 6216 7700
rect 6272 7672 6328 7700
rect 6356 7672 7084 7700
rect 6132 7644 6860 7672
rect 6888 7644 6972 7672
rect 5572 7616 5908 7644
rect 6104 7616 6748 7644
rect 6776 7616 6860 7644
rect 6916 7616 6972 7644
rect 7028 7644 7084 7672
rect 7140 7672 7196 7700
rect 7252 7672 7588 7700
rect 7644 7700 7700 7728
rect 7728 7700 7952 7728
rect 7644 7672 7952 7700
rect 8008 7700 8064 7728
rect 8092 7700 8316 7728
rect 8008 7672 8288 7700
rect 8344 7672 8568 7728
rect 8624 7700 8820 7728
rect 8876 7700 9352 7728
rect 8624 7672 8988 7700
rect 9016 7672 9352 7700
rect 7140 7644 7476 7672
rect 7532 7644 8204 7672
rect 8260 7644 8764 7672
rect 8820 7644 9352 7672
rect 9436 7700 9716 7728
rect 9436 7644 9744 7700
rect 9912 7644 9940 7700
rect 7028 7616 7364 7644
rect 1456 7588 2044 7616
rect 2268 7588 2464 7616
rect 3276 7588 3332 7616
rect 5432 7588 5880 7616
rect 1456 7560 2072 7588
rect 2324 7560 2352 7588
rect 2408 7560 2464 7588
rect 5376 7560 5516 7588
rect 1008 7532 1036 7560
rect 1204 7532 2072 7560
rect 2408 7532 2436 7560
rect 2660 7532 2688 7560
rect 5376 7532 5432 7560
rect 5460 7532 5516 7560
rect 5544 7532 5600 7588
rect 5628 7560 5880 7588
rect 5656 7532 5684 7560
rect 5740 7532 5768 7560
rect 5852 7532 5880 7560
rect 6076 7588 6272 7616
rect 6300 7588 6384 7616
rect 6076 7532 6132 7588
rect 6160 7532 6188 7588
rect 6244 7532 6272 7588
rect 6328 7560 6356 7588
rect 6412 7560 6524 7616
rect 6552 7588 6636 7616
rect 6664 7588 6748 7616
rect 6804 7588 6860 7616
rect 6888 7588 7252 7616
rect 6580 7560 6636 7588
rect 6692 7560 7140 7588
rect 7168 7560 7252 7588
rect 7308 7588 7364 7616
rect 7420 7616 7532 7644
rect 7616 7616 8232 7644
rect 8260 7616 8484 7644
rect 7420 7588 7504 7616
rect 7308 7560 7504 7588
rect 7644 7588 7756 7616
rect 7812 7588 8120 7616
rect 7644 7560 7672 7588
rect 7728 7560 8036 7588
rect 8064 7560 8120 7588
rect 8176 7588 8484 7616
rect 8512 7616 9772 7644
rect 8512 7588 8708 7616
rect 8764 7588 8932 7616
rect 8988 7588 9772 7616
rect 8176 7560 8400 7588
rect 8456 7560 8708 7588
rect 8736 7560 9800 7588
rect 6328 7532 6384 7560
rect 6412 7532 7000 7560
rect 7056 7532 7112 7560
rect 7196 7532 7532 7560
rect 7644 7532 8008 7560
rect 8064 7532 8316 7560
rect 8344 7532 8400 7560
rect 8428 7532 8652 7560
rect 8680 7532 8876 7560
rect 1176 7476 2072 7532
rect 2352 7476 2380 7504
rect 2632 7476 2716 7532
rect 5348 7504 5768 7532
rect 6076 7504 6888 7532
rect 5376 7476 5852 7504
rect 6104 7476 6300 7504
rect 6356 7476 6664 7504
rect 1176 7448 2044 7476
rect 2268 7448 2380 7476
rect 3976 7448 4004 7476
rect 4312 7448 4340 7476
rect 4872 7448 4928 7476
rect 5348 7448 5404 7476
rect 5460 7448 5488 7476
rect 1148 7420 2072 7448
rect 2240 7420 2380 7448
rect 5348 7420 5488 7448
rect 5544 7448 5600 7476
rect 5628 7448 5852 7476
rect 5544 7420 5684 7448
rect 5740 7420 5768 7448
rect 5824 7420 5880 7448
rect 6132 7420 6272 7476
rect 6356 7448 6384 7476
rect 6440 7420 6524 7476
rect 6608 7420 6664 7476
rect 6720 7448 6776 7504
rect 6832 7476 6888 7504
rect 6944 7504 7000 7532
rect 7084 7504 7532 7532
rect 7616 7504 7896 7532
rect 6944 7476 7420 7504
rect 7476 7476 7812 7504
rect 7840 7476 7896 7504
rect 7952 7504 8288 7532
rect 8372 7504 8876 7532
rect 8904 7532 9800 7560
rect 8904 7504 9828 7532
rect 7952 7476 8204 7504
rect 6832 7448 7280 7476
rect 7364 7448 7420 7476
rect 7448 7448 7784 7476
rect 6692 7420 7168 7448
rect 952 7392 1008 7420
rect 1148 7392 2044 7420
rect 2212 7392 2380 7420
rect 4088 7392 4116 7420
rect 5348 7392 5684 7420
rect 5712 7392 5796 7420
rect 5824 7392 5908 7420
rect 6412 7392 7056 7420
rect 1148 7364 1848 7392
rect 1988 7364 2044 7392
rect 1120 7336 1820 7364
rect 1960 7336 2044 7364
rect 2184 7336 2408 7392
rect 3696 7336 3752 7392
rect 5348 7364 5964 7392
rect 6384 7364 6832 7392
rect 6860 7364 6944 7392
rect 1120 7308 1792 7336
rect 1904 7308 2100 7336
rect 896 7280 924 7308
rect 1092 7280 1764 7308
rect 1092 7252 1736 7280
rect 1876 7252 2100 7308
rect 2240 7280 2408 7336
rect 5376 7308 5432 7364
rect 5488 7336 5544 7364
rect 5628 7336 5908 7364
rect 6244 7336 6580 7364
rect 6608 7336 6692 7364
rect 5488 7308 5516 7336
rect 5376 7280 5488 7308
rect 5656 7280 5684 7336
rect 5740 7280 5768 7336
rect 5796 7280 5880 7336
rect 6272 7280 6328 7336
rect 6384 7280 6440 7336
rect 6496 7308 6552 7336
rect 6636 7308 6692 7336
rect 6748 7308 6804 7364
rect 6888 7336 6944 7364
rect 7000 7364 7056 7392
rect 7112 7392 7168 7420
rect 7224 7420 7308 7448
rect 7336 7420 7672 7448
rect 7224 7392 7560 7420
rect 7112 7364 7476 7392
rect 7000 7336 7364 7364
rect 6860 7308 7224 7336
rect 6524 7280 6580 7308
rect 6608 7280 7112 7308
rect 7140 7280 7196 7308
rect 7280 7280 7336 7336
rect 7392 7308 7448 7364
rect 7504 7336 7560 7392
rect 7616 7392 7672 7420
rect 7728 7420 7784 7448
rect 7840 7448 8204 7476
rect 8260 7476 8316 7504
rect 8344 7476 8568 7504
rect 8260 7448 8596 7476
rect 8624 7448 8820 7504
rect 8848 7476 9044 7504
rect 9072 7476 9828 7504
rect 9912 7476 9968 7532
rect 8848 7448 9184 7476
rect 9212 7448 9828 7476
rect 7840 7420 8092 7448
rect 7728 7392 8008 7420
rect 8036 7392 8092 7420
rect 8148 7420 8484 7448
rect 8540 7420 8736 7448
rect 8148 7392 8400 7420
rect 8428 7392 8484 7420
rect 8512 7392 8736 7420
rect 8792 7392 8988 7448
rect 9016 7392 9856 7448
rect 7616 7364 7980 7392
rect 7616 7336 7868 7364
rect 7504 7308 7868 7336
rect 7924 7336 7980 7364
rect 8036 7364 8400 7392
rect 8456 7364 8680 7392
rect 8708 7364 9156 7392
rect 9184 7364 9884 7392
rect 10024 7364 10052 7392
rect 8036 7336 8288 7364
rect 7924 7308 8288 7336
rect 8344 7336 8652 7364
rect 8708 7336 8904 7364
rect 8960 7336 9884 7364
rect 8344 7308 8596 7336
rect 8624 7308 9072 7336
rect 9100 7308 9912 7336
rect 7392 7280 7728 7308
rect 2268 7252 2380 7280
rect 3192 7252 3248 7280
rect 3864 7252 3892 7280
rect 4452 7252 4480 7280
rect 4816 7252 4928 7280
rect 5376 7252 5460 7280
rect 5628 7252 5824 7280
rect 6244 7252 7000 7280
rect 1064 7224 1708 7252
rect 1876 7224 2044 7252
rect 2352 7224 2380 7252
rect 4816 7224 4900 7252
rect 1064 7196 1652 7224
rect 4788 7196 4900 7224
rect 5656 7224 5824 7252
rect 5656 7196 5712 7224
rect 5740 7196 5824 7224
rect 6188 7224 6720 7252
rect 6188 7196 6356 7224
rect 6384 7196 6468 7224
rect 1092 7168 1624 7196
rect 3360 7168 3388 7196
rect 4844 7168 4956 7196
rect 5656 7168 5684 7196
rect 504 7140 532 7168
rect 868 7140 896 7168
rect 1092 7140 1540 7168
rect 4844 7140 4928 7168
rect 5656 7140 5712 7168
rect 5740 7140 5796 7196
rect 6188 7168 6244 7196
rect 6272 7168 6328 7196
rect 6188 7140 6216 7168
rect 6300 7140 6328 7168
rect 6412 7140 6468 7196
rect 6524 7140 6580 7224
rect 6664 7168 6720 7224
rect 6776 7196 6832 7252
rect 6916 7196 6972 7252
rect 7028 7224 7084 7280
rect 7168 7252 7224 7280
rect 7280 7252 7616 7280
rect 7168 7224 7504 7252
rect 7560 7224 7616 7252
rect 7700 7252 7728 7280
rect 7812 7280 7868 7308
rect 7896 7280 8176 7308
rect 7812 7252 8176 7280
rect 8232 7280 8568 7308
rect 8624 7280 8848 7308
rect 8232 7252 8848 7280
rect 8876 7252 9912 7308
rect 7700 7224 8064 7252
rect 7028 7196 7392 7224
rect 7448 7196 7504 7224
rect 7588 7196 7644 7224
rect 7672 7196 7952 7224
rect 8008 7196 8064 7224
rect 8120 7224 8484 7252
rect 8540 7224 8764 7252
rect 8792 7224 9072 7252
rect 8120 7196 8372 7224
rect 8400 7196 8484 7224
rect 8512 7196 8764 7224
rect 8820 7196 9044 7224
rect 9128 7196 9548 7252
rect 9576 7224 9940 7252
rect 9604 7196 9940 7224
rect 6776 7168 6860 7196
rect 6888 7168 7280 7196
rect 7308 7168 7392 7196
rect 7476 7168 7504 7196
rect 7560 7168 7924 7196
rect 8008 7168 8372 7196
rect 8428 7168 8680 7196
rect 8708 7168 8904 7196
rect 8932 7168 9044 7196
rect 9100 7168 9968 7196
rect 6636 7140 7140 7168
rect 7196 7140 7252 7168
rect 1120 7112 1512 7140
rect 4172 7112 4228 7140
rect 4844 7112 4900 7140
rect 5516 7112 5544 7140
rect 5684 7112 5796 7140
rect 6160 7112 6244 7140
rect 6272 7112 6356 7140
rect 6384 7112 7028 7140
rect 812 7028 840 7084
rect 1008 7056 1064 7084
rect 1092 7056 1484 7112
rect 2296 7084 2324 7112
rect 2520 7056 2604 7084
rect 3528 7056 3556 7112
rect 4592 7056 4676 7084
rect 4872 7056 4900 7112
rect 5460 7084 5488 7112
rect 5684 7084 5768 7112
rect 6104 7084 6776 7112
rect 6804 7084 6860 7112
rect 1008 7028 1456 7056
rect 2492 7028 2604 7056
rect 1008 7000 1036 7028
rect 980 6944 1036 7000
rect 1120 7000 1456 7028
rect 2520 7000 2576 7028
rect 4564 7000 4704 7056
rect 4844 7028 4928 7056
rect 5432 7028 5488 7084
rect 5712 7056 5740 7084
rect 6132 7056 6244 7084
rect 6272 7056 6356 7084
rect 4872 7000 4956 7028
rect 5460 7000 5488 7028
rect 5628 7000 5656 7028
rect 6132 7000 6216 7056
rect 6272 7000 6328 7056
rect 6412 7000 6468 7084
rect 6552 7000 6608 7084
rect 6692 7056 6720 7084
rect 6832 7056 6860 7084
rect 6944 7056 7000 7112
rect 7084 7084 7140 7140
rect 7224 7112 7252 7140
rect 7336 7140 7392 7168
rect 7448 7140 7812 7168
rect 7336 7112 7700 7140
rect 7196 7084 7588 7112
rect 7616 7084 7700 7112
rect 7756 7112 7812 7140
rect 7868 7140 7952 7168
rect 7980 7140 8260 7168
rect 7868 7112 8260 7140
rect 8316 7140 8652 7168
rect 8708 7140 9968 7168
rect 8316 7112 8568 7140
rect 8596 7112 9968 7140
rect 7756 7084 8148 7112
rect 8204 7084 8568 7112
rect 8624 7084 9016 7112
rect 9044 7084 9996 7112
rect 7084 7056 7448 7084
rect 6692 7028 6748 7056
rect 6832 7028 6888 7056
rect 6944 7028 7336 7056
rect 7364 7028 7420 7056
rect 7504 7028 7560 7084
rect 7644 7056 8036 7084
rect 8064 7056 8148 7084
rect 8176 7056 8456 7084
rect 8484 7056 9996 7084
rect 7616 7028 8008 7056
rect 8064 7028 8456 7056
rect 8512 7028 8960 7056
rect 8988 7028 9156 7056
rect 9184 7028 9996 7056
rect 10136 7028 10192 7056
rect 6664 7000 7168 7028
rect 1120 6944 1428 7000
rect 1708 6944 1736 7000
rect 4564 6972 4676 7000
rect 2212 6944 2268 6972
rect 4592 6944 4648 6972
rect 4900 6944 4956 7000
rect 6132 6972 7056 7000
rect 6104 6944 6776 6972
rect 6832 6944 6916 6972
rect 980 6916 1008 6944
rect 952 6888 1008 6916
rect 1120 6916 1372 6944
rect 2184 6916 2296 6944
rect 1120 6888 1344 6916
rect 2212 6888 2268 6916
rect 2744 6888 2772 6944
rect 3892 6888 3920 6944
rect 4564 6916 4648 6944
rect 4872 6916 4956 6944
rect 5488 6916 5516 6944
rect 6076 6916 6132 6944
rect 6160 6916 6496 6944
rect 6580 6916 6636 6944
rect 6692 6916 6748 6944
rect 6860 6916 6888 6944
rect 6972 6916 7028 6972
rect 7112 6944 7168 7000
rect 7252 6972 7308 7028
rect 7392 7000 7448 7028
rect 7504 7000 7896 7028
rect 7364 6972 7756 7000
rect 7252 6944 7644 6972
rect 7672 6944 7756 6972
rect 7812 6972 7896 7000
rect 7924 7000 8344 7028
rect 8372 7000 8456 7028
rect 8484 7000 8736 7028
rect 8820 7000 8848 7028
rect 8876 7000 10024 7028
rect 7924 6972 8316 7000
rect 8372 6972 8736 7000
rect 8904 6972 9156 7000
rect 9240 6972 10024 7000
rect 7812 6944 8204 6972
rect 7112 6916 7504 6944
rect 7532 6916 7616 6944
rect 7672 6916 8092 6944
rect 8120 6916 8204 6944
rect 8260 6944 8344 6972
rect 8372 6944 8624 6972
rect 8260 6916 8624 6944
rect 4508 6888 4620 6916
rect 4760 6888 4816 6916
rect 4844 6888 4984 6916
rect 5460 6888 5544 6916
rect 5628 6888 5684 6916
rect 5824 6888 5852 6916
rect 756 6832 812 6888
rect 952 6832 980 6888
rect 1148 6860 1344 6888
rect 4508 6860 4564 6888
rect 1148 6832 1316 6860
rect 4088 6832 4116 6860
rect 4760 6832 4844 6888
rect 4872 6860 4984 6888
rect 5432 6860 5712 6888
rect 5768 6860 5852 6888
rect 5908 6888 5964 6916
rect 5908 6860 5992 6888
rect 6076 6860 6104 6916
rect 6188 6860 6216 6916
rect 6300 6860 6356 6916
rect 6440 6888 6468 6916
rect 6580 6888 6608 6916
rect 6720 6888 6748 6916
rect 6832 6888 6916 6916
rect 6972 6888 7364 6916
rect 6440 6860 6496 6888
rect 6552 6860 6636 6888
rect 6692 6860 7224 6888
rect 7280 6860 7336 6888
rect 7420 6860 7504 6916
rect 7560 6888 7644 6916
rect 7672 6888 8064 6916
rect 8148 6888 8512 6916
rect 7532 6860 7952 6888
rect 4872 6832 5012 6860
rect 5432 6832 6244 6860
rect 6272 6832 6384 6860
rect 6412 6832 7084 6860
rect 924 6748 952 6832
rect 1148 6804 1260 6832
rect 2408 6804 2464 6832
rect 4760 6804 5012 6832
rect 5292 6804 5348 6832
rect 5432 6804 5460 6832
rect 5544 6804 5572 6832
rect 1148 6776 1232 6804
rect 3416 6776 3444 6804
rect 896 6720 952 6748
rect 728 6664 756 6692
rect 896 6636 924 6720
rect 868 6580 924 6636
rect 1120 6692 1204 6776
rect 1904 6748 1932 6776
rect 4760 6748 4956 6804
rect 5292 6776 5376 6804
rect 5404 6776 5460 6804
rect 5516 6776 5572 6804
rect 5628 6804 5684 6832
rect 5628 6776 5656 6804
rect 5712 6776 5768 6832
rect 5824 6804 6804 6832
rect 6860 6804 6944 6832
rect 5852 6776 5880 6804
rect 5236 6748 5768 6776
rect 5824 6748 5880 6776
rect 5936 6748 5992 6804
rect 6076 6776 6132 6804
rect 6188 6776 6244 6804
rect 6300 6776 6384 6804
rect 6440 6776 6524 6804
rect 6076 6748 6104 6776
rect 6188 6748 6216 6776
rect 6300 6748 6356 6776
rect 4760 6720 4788 6748
rect 4844 6720 5012 6748
rect 5208 6720 5236 6748
rect 3108 6692 3136 6720
rect 4844 6692 4984 6720
rect 5124 6692 5236 6720
rect 5292 6720 5348 6748
rect 5376 6720 5992 6748
rect 6048 6720 6132 6748
rect 6188 6720 6244 6748
rect 6300 6720 6384 6748
rect 6440 6720 6496 6776
rect 6580 6720 6664 6804
rect 6720 6776 6776 6804
rect 6888 6776 6944 6804
rect 7028 6776 7084 6832
rect 7140 6832 7196 6860
rect 7280 6832 7364 6860
rect 7392 6832 7812 6860
rect 7140 6804 7224 6832
rect 7280 6804 7700 6832
rect 7728 6804 7812 6832
rect 7868 6832 7952 6860
rect 8008 6860 8092 6888
rect 8120 6860 8512 6888
rect 8568 6888 8624 6916
rect 8680 6944 8736 6972
rect 8820 6944 8848 6972
rect 8876 6944 9128 6972
rect 9240 6944 10052 6972
rect 8680 6916 9128 6944
rect 8680 6888 8988 6916
rect 8568 6860 8988 6888
rect 9016 6888 9156 6916
rect 9212 6888 10052 6944
rect 9016 6860 9184 6888
rect 9212 6860 10080 6888
rect 8008 6832 8400 6860
rect 7868 6804 8288 6832
rect 8316 6804 8400 6832
rect 8456 6832 8904 6860
rect 8932 6832 9100 6860
rect 9128 6832 10080 6860
rect 8456 6804 8792 6832
rect 7140 6776 7560 6804
rect 7588 6776 7672 6804
rect 6748 6748 6804 6776
rect 6860 6748 7420 6776
rect 7448 6748 7532 6776
rect 7616 6748 7672 6776
rect 7728 6776 8288 6804
rect 8344 6776 8792 6804
rect 8848 6776 10080 6832
rect 7728 6748 8148 6776
rect 6720 6720 7280 6748
rect 7336 6720 7392 6748
rect 7476 6720 7560 6748
rect 7588 6720 8148 6748
rect 8204 6748 8288 6776
rect 8316 6748 8708 6776
rect 8764 6748 9044 6776
rect 9072 6748 9128 6776
rect 9156 6748 9352 6776
rect 9380 6748 10108 6776
rect 10220 6748 10276 6804
rect 8204 6720 8596 6748
rect 5292 6692 5320 6720
rect 1120 6636 1176 6692
rect 1988 6636 2016 6692
rect 5096 6664 5320 6692
rect 5404 6692 5460 6720
rect 5488 6692 7112 6720
rect 5404 6664 5432 6692
rect 5516 6664 5628 6692
rect 5684 6664 5768 6692
rect 1120 6580 1204 6636
rect 3780 6608 3836 6664
rect 5068 6636 5460 6664
rect 5488 6636 5768 6664
rect 5824 6664 5908 6692
rect 5964 6664 6048 6692
rect 6076 6664 6860 6692
rect 5824 6636 5880 6664
rect 5040 6608 5152 6636
rect 5208 6608 5908 6636
rect 5964 6608 6020 6664
rect 6104 6636 6160 6664
rect 6188 6636 6272 6664
rect 6104 6608 6132 6636
rect 6216 6608 6244 6636
rect 3332 6580 3360 6608
rect 868 6552 896 6580
rect 1148 6552 1176 6580
rect 5012 6552 5152 6608
rect 5236 6580 5264 6608
rect 5208 6552 5264 6580
rect 5348 6580 5404 6608
rect 5460 6580 6160 6608
rect 6188 6580 6272 6608
rect 6328 6580 6384 6664
rect 6468 6636 6552 6664
rect 6608 6636 6692 6664
rect 6468 6580 6524 6636
rect 6636 6608 6664 6636
rect 6776 6608 6832 6664
rect 6916 6608 6972 6692
rect 7056 6636 7112 6692
rect 7196 6692 7252 6720
rect 7336 6692 7420 6720
rect 7448 6692 8036 6720
rect 8092 6692 8596 6720
rect 8652 6720 8708 6748
rect 8736 6720 9044 6748
rect 9100 6720 10108 6748
rect 8652 6692 8960 6720
rect 7196 6664 7280 6692
rect 7336 6664 7728 6692
rect 7168 6636 7616 6664
rect 7028 6608 7588 6636
rect 6608 6580 6692 6608
rect 6748 6580 7336 6608
rect 5348 6552 5376 6580
rect 840 6440 896 6552
rect 1120 6496 1176 6552
rect 1428 6496 1540 6552
rect 2492 6524 2520 6552
rect 4956 6524 5292 6552
rect 5320 6524 5376 6552
rect 5460 6524 5516 6580
rect 1428 6440 1512 6496
rect 2464 6468 2548 6524
rect 2996 6496 3052 6524
rect 4816 6496 5012 6524
rect 4228 6468 4256 6496
rect 4704 6468 5012 6496
rect 5068 6496 5544 6524
rect 5572 6496 5628 6580
rect 5684 6552 5740 6580
rect 5824 6552 6552 6580
rect 6580 6552 7168 6580
rect 5712 6524 5740 6552
rect 5684 6496 5740 6524
rect 5852 6496 5908 6552
rect 5936 6524 6888 6552
rect 6916 6524 7028 6552
rect 5964 6496 6020 6524
rect 5068 6468 5124 6496
rect 2492 6440 2520 6468
rect 2716 6440 2744 6468
rect 4732 6440 5124 6468
rect 5180 6468 5264 6496
rect 5292 6468 5404 6496
rect 5432 6468 5740 6496
rect 5824 6468 6020 6496
rect 6076 6468 6160 6524
rect 5180 6440 5236 6468
rect 840 6328 868 6440
rect 924 6412 952 6440
rect 2660 6412 2772 6440
rect 3668 6412 3752 6440
rect 4788 6412 5236 6440
rect 5320 6412 5348 6468
rect 924 6328 980 6412
rect 2632 6384 2772 6412
rect 672 6272 700 6300
rect 896 6272 980 6328
rect 2604 6328 2660 6384
rect 2716 6328 2772 6384
rect 3416 6328 3472 6356
rect 3640 6328 3780 6412
rect 4816 6384 5376 6412
rect 5460 6384 5488 6468
rect 5572 6440 5656 6468
rect 5684 6440 6160 6468
rect 6216 6468 6300 6524
rect 6356 6496 6440 6524
rect 6496 6496 6580 6524
rect 6636 6496 6720 6524
rect 6776 6496 6860 6524
rect 6356 6468 6412 6496
rect 6216 6440 6412 6468
rect 6496 6440 6552 6496
rect 6664 6468 6720 6496
rect 6804 6468 6860 6496
rect 6944 6496 7000 6524
rect 7084 6496 7168 6552
rect 7224 6524 7308 6580
rect 7364 6552 7448 6608
rect 7504 6580 7588 6608
rect 7644 6608 7728 6664
rect 7784 6664 7896 6692
rect 7924 6664 8036 6692
rect 8064 6664 8484 6692
rect 7784 6636 8372 6664
rect 8400 6636 8484 6664
rect 8540 6664 8596 6692
rect 8624 6664 8960 6692
rect 9016 6692 9464 6720
rect 9492 6692 10108 6720
rect 9016 6664 9296 6692
rect 9324 6664 10108 6692
rect 10248 6664 10276 6692
rect 8540 6636 8876 6664
rect 8932 6636 9212 6664
rect 7756 6608 8344 6636
rect 8428 6608 8792 6636
rect 8820 6608 8876 6636
rect 8904 6608 9212 6636
rect 9240 6636 10136 6664
rect 9240 6608 9408 6636
rect 9436 6608 10136 6636
rect 7644 6580 8232 6608
rect 7504 6552 8120 6580
rect 8148 6552 8232 6580
rect 8288 6580 8344 6608
rect 8400 6580 8764 6608
rect 8820 6580 9128 6608
rect 8288 6552 8652 6580
rect 8736 6552 9044 6580
rect 7364 6524 7896 6552
rect 7224 6496 7784 6524
rect 7952 6496 8092 6552
rect 8176 6524 8568 6552
rect 8596 6524 8652 6552
rect 8708 6524 9044 6552
rect 9072 6552 9128 6580
rect 9156 6580 10136 6608
rect 9156 6552 9352 6580
rect 9380 6552 10136 6580
rect 9072 6524 10164 6552
rect 8148 6496 8540 6524
rect 8624 6496 8932 6524
rect 6944 6468 7028 6496
rect 7084 6468 7644 6496
rect 6636 6440 6720 6468
rect 6776 6440 7644 6468
rect 7672 6468 7784 6496
rect 8036 6468 8428 6496
rect 7672 6440 7728 6468
rect 8036 6440 8316 6468
rect 8344 6440 8428 6468
rect 8484 6468 8540 6496
rect 8596 6468 8932 6496
rect 8988 6468 9268 6524
rect 9296 6468 10164 6524
rect 8484 6440 8848 6468
rect 8904 6440 9184 6468
rect 5572 6384 5628 6440
rect 5712 6412 7280 6440
rect 7308 6412 7392 6440
rect 7448 6412 7728 6440
rect 8064 6412 8176 6440
rect 8204 6412 8288 6440
rect 8372 6412 8428 6440
rect 8456 6412 8736 6440
rect 5684 6384 5880 6412
rect 5936 6384 7700 6412
rect 4536 6356 4564 6384
rect 4816 6328 4872 6384
rect 4928 6356 4984 6384
rect 4900 6328 4984 6356
rect 5068 6356 7028 6384
rect 7084 6356 7672 6384
rect 8092 6356 8148 6412
rect 8232 6384 8288 6412
rect 8344 6384 8736 6412
rect 8792 6412 8848 6440
rect 8876 6412 9184 6440
rect 9212 6440 10164 6468
rect 9212 6412 9380 6440
rect 9408 6412 10164 6440
rect 8792 6384 9100 6412
rect 8232 6356 8624 6384
rect 5068 6328 5124 6356
rect 5180 6328 5236 6356
rect 2604 6300 2772 6328
rect 3668 6300 3752 6328
rect 2632 6272 2744 6300
rect 3892 6272 3948 6328
rect 4788 6300 5012 6328
rect 5040 6300 5124 6328
rect 5152 6300 5236 6328
rect 5292 6328 6720 6356
rect 5292 6300 5376 6328
rect 4788 6272 5376 6300
rect 5432 6272 5488 6328
rect 5572 6300 5740 6328
rect 5572 6272 5628 6300
rect 868 6244 980 6272
rect 840 6216 980 6244
rect 2072 6216 2128 6272
rect 4788 6216 4844 6272
rect 4900 6244 5208 6272
rect 5264 6244 5628 6272
rect 5684 6244 5740 6300
rect 5824 6300 5908 6328
rect 5936 6300 5992 6328
rect 6076 6300 6300 6328
rect 5824 6244 5852 6300
rect 4900 6216 4956 6244
rect 644 6132 672 6160
rect 840 6132 952 6216
rect 3164 6160 3192 6188
rect 4200 6160 4228 6216
rect 4788 6188 4956 6216
rect 5012 6188 5096 6244
rect 5124 6188 5180 6244
rect 4368 6160 4424 6188
rect 616 5880 672 5908
rect 868 5880 952 6132
rect 1092 6104 1120 6160
rect 1064 6076 1148 6104
rect 2324 6076 2352 6104
rect 2828 6076 2884 6160
rect 4340 6132 4508 6160
rect 4760 6132 5180 6188
rect 5292 6216 5768 6244
rect 5796 6216 5880 6244
rect 5964 6216 5992 6300
rect 6104 6244 6160 6300
rect 6244 6272 6300 6300
rect 6216 6244 6300 6272
rect 6356 6244 6440 6328
rect 6524 6272 6608 6328
rect 6636 6300 6720 6328
rect 6804 6328 6888 6356
rect 6916 6328 7056 6356
rect 7084 6328 7616 6356
rect 8092 6328 8176 6356
rect 8204 6328 8512 6356
rect 8540 6328 8624 6356
rect 8680 6356 8736 6384
rect 8764 6356 9016 6384
rect 9044 6356 9100 6384
rect 9128 6384 10164 6412
rect 9128 6356 9296 6384
rect 9352 6356 10192 6384
rect 8680 6328 8988 6356
rect 9044 6328 9492 6356
rect 9520 6328 10192 6356
rect 6804 6300 6944 6328
rect 6636 6272 6748 6300
rect 6776 6272 6944 6300
rect 7028 6300 7420 6328
rect 7448 6300 7588 6328
rect 8092 6300 8484 6328
rect 8568 6300 8904 6328
rect 7028 6272 7252 6300
rect 7336 6272 7392 6300
rect 6524 6244 6664 6272
rect 6720 6244 6888 6272
rect 7084 6244 7252 6272
rect 7308 6244 7392 6272
rect 7476 6244 7560 6300
rect 7924 6272 8008 6300
rect 8064 6272 8372 6300
rect 8428 6272 8484 6300
rect 8540 6272 8904 6300
rect 8960 6272 9240 6328
rect 9268 6300 10192 6328
rect 9268 6272 10164 6300
rect 7924 6244 8232 6272
rect 6104 6216 6636 6244
rect 6776 6216 6832 6244
rect 7084 6216 7588 6244
rect 7924 6216 8092 6244
rect 8148 6216 8232 6244
rect 5292 6188 6608 6216
rect 6804 6188 6832 6216
rect 7056 6188 7588 6216
rect 5292 6160 5572 6188
rect 5712 6160 6440 6188
rect 5292 6132 5544 6160
rect 5712 6132 5852 6160
rect 5908 6132 5964 6160
rect 6020 6132 6104 6160
rect 6160 6132 6216 6160
rect 6272 6132 6328 6160
rect 6384 6132 6440 6160
rect 6524 6160 6580 6188
rect 6776 6160 6832 6188
rect 7000 6160 7588 6188
rect 7728 6160 7756 6216
rect 7952 6188 8092 6216
rect 8176 6188 8232 6216
rect 8288 6244 8344 6272
rect 8428 6244 8792 6272
rect 8288 6188 8680 6244
rect 7980 6160 8092 6188
rect 8148 6160 8568 6188
rect 8624 6160 8680 6188
rect 8736 6216 8792 6244
rect 8848 6244 9156 6272
rect 9184 6244 10164 6272
rect 8848 6216 9352 6244
rect 9380 6216 10136 6244
rect 8736 6188 9044 6216
rect 9100 6188 10164 6216
rect 10360 6188 10388 6244
rect 8736 6160 8960 6188
rect 8988 6160 9044 6188
rect 9072 6160 9268 6188
rect 9324 6160 10136 6188
rect 6524 6132 6552 6160
rect 6776 6132 6860 6160
rect 7000 6132 7336 6160
rect 4340 6104 4620 6132
rect 4732 6104 4844 6132
rect 4340 6076 4368 6104
rect 4424 6076 4816 6104
rect 4872 6076 4956 6132
rect 4984 6104 5236 6132
rect 5264 6104 5348 6132
rect 5404 6104 5544 6132
rect 5684 6104 6104 6132
rect 6132 6104 6468 6132
rect 6496 6104 6524 6132
rect 6804 6104 6832 6132
rect 7084 6104 7168 6132
rect 7252 6104 7308 6132
rect 5012 6076 5068 6104
rect 5096 6076 5320 6104
rect 5432 6076 5544 6104
rect 5740 6076 6524 6104
rect 6580 6076 6608 6104
rect 7252 6076 7280 6104
rect 7364 6076 7448 6160
rect 7504 6132 7616 6160
rect 8008 6132 8428 6160
rect 7504 6104 7644 6132
rect 8064 6104 8288 6132
rect 7504 6076 7672 6104
rect 8092 6076 8148 6104
rect 8204 6076 8288 6104
rect 1036 6048 1148 6076
rect 1876 6048 1904 6076
rect 4340 6048 4396 6076
rect 4424 6048 4452 6076
rect 4536 6048 4956 6076
rect 4984 6048 5040 6076
rect 5124 6048 5236 6076
rect 1036 6020 1176 6048
rect 1036 5992 1148 6020
rect 1848 5992 1932 6048
rect 3108 6020 3136 6048
rect 3612 6020 3668 6048
rect 4340 6020 4452 6048
rect 4508 6020 4564 6048
rect 3080 5992 3164 6020
rect 3808 5992 3836 6020
rect 1064 5964 1120 5992
rect 1512 5964 1540 5992
rect 2520 5936 2604 5992
rect 3080 5964 3136 5992
rect 4312 5964 4564 6020
rect 4620 6020 4984 6048
rect 5152 6020 5236 6048
rect 5432 6048 5572 6076
rect 5740 6048 6468 6076
rect 7252 6048 7700 6076
rect 5432 6020 5460 6048
rect 5488 6020 5572 6048
rect 4620 5964 4676 6020
rect 4732 5992 4984 6020
rect 5460 5992 5572 6020
rect 5852 6020 6328 6048
rect 6384 6020 6468 6048
rect 7224 6020 7728 6048
rect 8092 6020 8120 6076
rect 8232 6048 8288 6076
rect 8344 6076 8428 6132
rect 8484 6132 8540 6160
rect 8624 6132 8960 6160
rect 9016 6132 9492 6160
rect 9520 6132 10136 6160
rect 8484 6076 8848 6132
rect 8904 6104 8960 6132
rect 8988 6104 9184 6132
rect 9240 6104 10108 6132
rect 8904 6076 9212 6104
rect 9240 6076 9408 6104
rect 9436 6076 9576 6104
rect 9604 6076 10108 6104
rect 8344 6048 8736 6076
rect 8204 6020 8624 6048
rect 8652 6020 8736 6048
rect 8792 6048 8848 6076
rect 8876 6048 9100 6076
rect 9156 6048 10108 6076
rect 8792 6020 9100 6048
rect 9128 6020 9324 6048
rect 9352 6020 10080 6048
rect 5852 5992 5936 6020
rect 5992 5992 6104 6020
rect 6160 5992 6216 6020
rect 6272 5992 6328 6020
rect 6412 5992 6468 6020
rect 4732 5964 4816 5992
rect 3976 5936 4004 5964
rect 4284 5936 4340 5964
rect 2520 5908 2576 5936
rect 1008 5880 1036 5908
rect 4116 5880 4172 5936
rect 4256 5908 4340 5936
rect 4396 5936 4816 5964
rect 4844 5936 4900 5992
rect 5460 5964 5628 5992
rect 5824 5964 6328 5992
rect 6384 5964 6468 5992
rect 5488 5936 5628 5964
rect 5852 5936 6468 5964
rect 4396 5908 4424 5936
rect 4256 5880 4424 5908
rect 4480 5908 4956 5936
rect 5488 5908 5516 5936
rect 5572 5908 5628 5936
rect 5936 5908 6468 5936
rect 7308 5992 7756 6020
rect 8036 5992 8148 6020
rect 8176 5992 8596 6020
rect 8680 5992 8988 6020
rect 7308 5936 7364 5992
rect 7420 5936 7476 5992
rect 7560 5964 7616 5992
rect 7644 5964 7812 5992
rect 8036 5964 8064 5992
rect 8120 5964 8456 5992
rect 8540 5964 8596 5992
rect 8652 5964 8988 5992
rect 9044 5992 10108 6020
rect 9044 5964 9240 5992
rect 9296 5964 9464 5992
rect 7532 5936 7840 5964
rect 7308 5908 7840 5936
rect 8148 5936 8344 5964
rect 4480 5880 4536 5908
rect 616 5852 644 5880
rect 896 5852 1064 5880
rect 4256 5852 4536 5880
rect 4592 5880 4872 5908
rect 5348 5880 5404 5908
rect 5572 5880 5656 5908
rect 5964 5880 5992 5908
rect 6048 5880 6244 5908
rect 6272 5880 6356 5908
rect 4592 5852 4648 5880
rect 560 5740 588 5796
rect 896 5768 952 5852
rect 1008 5824 1064 5852
rect 2212 5824 2268 5852
rect 4256 5824 4312 5852
rect 4340 5824 4648 5852
rect 4704 5852 4788 5880
rect 5348 5852 5376 5880
rect 5600 5852 5656 5880
rect 4704 5824 4760 5852
rect 2212 5796 2240 5824
rect 2744 5768 2800 5824
rect 896 5740 980 5768
rect 2996 5740 3080 5824
rect 3164 5768 3248 5824
rect 4256 5796 4284 5824
rect 4340 5796 4396 5824
rect 4256 5768 4396 5796
rect 4452 5768 4760 5824
rect 5096 5796 5152 5852
rect 5320 5824 5376 5852
rect 5656 5824 5712 5852
rect 6048 5824 6104 5880
rect 6160 5824 6216 5880
rect 6272 5852 6328 5880
rect 6244 5824 6328 5852
rect 6384 5824 6468 5908
rect 7280 5880 7868 5908
rect 6832 5852 7028 5880
rect 7252 5852 7784 5880
rect 6748 5824 7532 5852
rect 7560 5824 7644 5852
rect 5292 5796 5404 5824
rect 5320 5768 5404 5796
rect 5600 5796 5740 5824
rect 6020 5796 6496 5824
rect 6580 5796 6664 5824
rect 6720 5796 7084 5824
rect 7112 5796 7392 5824
rect 5600 5768 5768 5796
rect 6020 5768 6328 5796
rect 6356 5768 6496 5796
rect 6720 5768 6804 5796
rect 6860 5768 6944 5796
rect 3192 5740 3220 5768
rect 4256 5740 4480 5768
rect 4536 5740 4732 5768
rect 588 5628 644 5656
rect 924 5628 952 5740
rect 2464 5712 2492 5740
rect 2996 5712 3052 5740
rect 3696 5712 3752 5740
rect 4340 5712 4620 5740
rect 4648 5712 4704 5740
rect 4872 5712 4900 5740
rect 5320 5712 5376 5768
rect 5656 5740 5852 5768
rect 6020 5740 6300 5768
rect 6440 5740 6468 5768
rect 6748 5740 6776 5768
rect 5684 5712 5796 5740
rect 4340 5684 4368 5712
rect 1148 5656 1176 5684
rect 4424 5656 4676 5712
rect 4844 5656 4928 5712
rect 5292 5684 5320 5712
rect 5348 5684 5376 5712
rect 5712 5684 5796 5712
rect 6020 5684 6188 5740
rect 6720 5712 6776 5740
rect 6860 5740 6916 5768
rect 7000 5740 7056 5796
rect 7140 5768 7224 5796
rect 7280 5768 7392 5796
rect 7448 5796 7504 5824
rect 7588 5796 7644 5824
rect 7728 5824 7784 5852
rect 8148 5852 8204 5936
rect 8260 5908 8344 5936
rect 8400 5936 8484 5964
rect 8540 5936 8876 5964
rect 8400 5908 8792 5936
rect 8820 5908 8876 5936
rect 8932 5936 9464 5964
rect 9492 5936 10108 5992
rect 10360 5936 10416 5964
rect 8932 5908 9128 5936
rect 9184 5908 9380 5936
rect 8288 5880 8344 5908
rect 8372 5880 8764 5908
rect 8260 5852 8652 5880
rect 8148 5824 8540 5852
rect 7728 5796 7812 5824
rect 7448 5768 7532 5796
rect 7560 5768 7644 5796
rect 7700 5768 7812 5796
rect 8176 5796 8400 5824
rect 8428 5796 8512 5824
rect 8176 5768 8260 5796
rect 7140 5740 7812 5768
rect 8204 5740 8232 5768
rect 6860 5712 6944 5740
rect 6972 5712 7868 5740
rect 8176 5712 8232 5740
rect 8316 5740 8372 5796
rect 8456 5768 8512 5796
rect 8568 5796 8652 5852
rect 8708 5852 8764 5880
rect 8820 5880 9380 5908
rect 9408 5908 10108 5936
rect 9408 5880 9576 5908
rect 9604 5880 10136 5908
rect 10192 5880 10220 5908
rect 8820 5852 9044 5880
rect 8708 5824 9016 5852
rect 9072 5824 9296 5880
rect 9324 5852 10136 5880
rect 10164 5852 10220 5880
rect 9324 5824 9492 5852
rect 9548 5824 10164 5852
rect 10192 5824 10220 5852
rect 8680 5796 8932 5824
rect 8568 5768 8932 5796
rect 8988 5796 9044 5824
rect 9072 5796 9212 5824
rect 8988 5768 9212 5796
rect 9240 5796 10136 5824
rect 9240 5768 9436 5796
rect 8456 5740 8820 5768
rect 8848 5740 8932 5768
rect 8960 5740 9100 5768
rect 9156 5740 9436 5768
rect 9464 5768 9968 5796
rect 9996 5768 10136 5796
rect 9464 5740 9940 5768
rect 8316 5712 8792 5740
rect 8876 5712 9072 5740
rect 6468 5684 7840 5712
rect 8176 5684 8680 5712
rect 1820 5628 1848 5656
rect 4060 5628 4088 5656
rect 4368 5628 4452 5656
rect 4508 5628 4536 5656
rect 588 5600 616 5628
rect 868 5488 952 5628
rect 2688 5600 2716 5628
rect 1372 5572 1400 5600
rect 5740 5572 5796 5684
rect 5992 5656 6216 5684
rect 6104 5600 6216 5656
rect 6076 5572 6216 5600
rect 6468 5656 7420 5684
rect 6468 5600 7084 5656
rect 7168 5628 7308 5656
rect 7364 5628 7420 5656
rect 7504 5628 7560 5684
rect 7616 5656 7812 5684
rect 8148 5656 8568 5684
rect 8596 5656 8680 5684
rect 8736 5684 8820 5712
rect 8848 5684 9072 5712
rect 8736 5656 9072 5684
rect 9156 5656 9912 5740
rect 10024 5712 10136 5768
rect 10080 5656 10136 5712
rect 7644 5628 7812 5656
rect 7896 5628 7952 5656
rect 8092 5628 8428 5656
rect 8456 5628 8540 5656
rect 8624 5628 8960 5656
rect 7168 5600 7448 5628
rect 7476 5600 7560 5628
rect 7616 5600 8008 5628
rect 8064 5600 8288 5628
rect 8316 5600 8400 5628
rect 6468 5572 6524 5600
rect 4228 5544 4256 5572
rect 5628 5544 5656 5572
rect 868 5460 924 5488
rect 2940 5460 2968 5488
rect 3472 5460 3528 5544
rect 4396 5516 4452 5544
rect 4564 5516 4620 5544
rect 5600 5516 5712 5544
rect 6104 5516 6244 5572
rect 6496 5544 6524 5572
rect 6580 5544 6664 5600
rect 6692 5572 7000 5600
rect 7028 5572 7112 5600
rect 7140 5572 8148 5600
rect 8176 5572 8260 5600
rect 6720 5544 8008 5572
rect 6524 5516 7728 5544
rect 3640 5488 3668 5516
rect 3864 5488 3920 5516
rect 4368 5488 4480 5516
rect 4536 5488 4620 5516
rect 4704 5488 5068 5516
rect 5096 5488 5236 5516
rect 5628 5488 5712 5516
rect 5964 5488 5992 5516
rect 6104 5488 6188 5516
rect 6216 5488 6244 5516
rect 6328 5488 6412 5516
rect 588 5432 644 5460
rect 588 5404 616 5432
rect 1428 5404 1456 5460
rect 3836 5432 3948 5488
rect 4368 5460 5264 5488
rect 5320 5460 5376 5488
rect 6104 5460 6132 5488
rect 6160 5460 6188 5488
rect 6356 5460 6412 5488
rect 6524 5488 7000 5516
rect 7084 5488 7308 5516
rect 7364 5488 7448 5516
rect 6524 5460 6748 5488
rect 6804 5460 6916 5488
rect 7140 5460 7196 5488
rect 7252 5460 7308 5488
rect 7392 5460 7448 5488
rect 7532 5460 7588 5516
rect 7672 5460 7728 5516
rect 7784 5488 7868 5544
rect 7924 5488 7980 5544
rect 8064 5516 8120 5572
rect 8204 5544 8260 5572
rect 8344 5572 8400 5600
rect 8484 5600 8568 5628
rect 8596 5600 8960 5628
rect 9016 5628 9100 5656
rect 9128 5628 9352 5656
rect 9436 5628 9464 5656
rect 9492 5628 9632 5656
rect 9660 5628 9856 5656
rect 9016 5600 9184 5628
rect 9212 5600 9352 5628
rect 9464 5600 9856 5628
rect 10080 5628 10164 5656
rect 10080 5600 10220 5628
rect 8484 5572 8848 5600
rect 8344 5544 8736 5572
rect 8764 5544 8848 5572
rect 8904 5544 9380 5600
rect 9464 5572 9744 5600
rect 9772 5572 9828 5600
rect 9436 5544 9576 5572
rect 9604 5544 9828 5572
rect 8204 5516 8708 5544
rect 8792 5516 9100 5544
rect 8064 5488 8596 5516
rect 7784 5460 8456 5488
rect 4340 5432 5376 5460
rect 6524 5432 6608 5460
rect 6832 5432 6860 5460
rect 7168 5432 7336 5460
rect 7364 5432 8344 5460
rect 3836 5404 3920 5432
rect 4312 5404 4396 5432
rect 1400 5376 1456 5404
rect 4256 5376 4396 5404
rect 2604 5348 2632 5376
rect 4228 5348 4396 5376
rect 4480 5404 5376 5432
rect 7140 5404 8204 5432
rect 4480 5376 4564 5404
rect 4592 5376 5404 5404
rect 4480 5348 4536 5376
rect 4592 5348 4676 5376
rect 4200 5320 4676 5348
rect 4732 5348 5404 5376
rect 7140 5376 7924 5404
rect 7140 5348 7504 5376
rect 7532 5348 7644 5376
rect 7672 5348 7756 5376
rect 4732 5320 4816 5348
rect 616 5292 644 5320
rect 980 5292 1008 5320
rect 952 5264 1036 5292
rect 952 5236 1064 5264
rect 1400 5236 1456 5320
rect 3192 5292 3220 5320
rect 4200 5292 4816 5320
rect 4844 5292 4900 5348
rect 2856 5236 2884 5264
rect 3388 5236 3444 5292
rect 4004 5264 4032 5292
rect 4116 5264 4144 5292
rect 4228 5264 4900 5292
rect 4984 5320 5320 5348
rect 5656 5320 5684 5348
rect 6244 5320 6356 5348
rect 6496 5320 6524 5348
rect 6860 5320 6972 5348
rect 7196 5320 7364 5348
rect 4984 5264 5152 5320
rect 4116 5236 4172 5264
rect 4228 5236 4312 5264
rect 4340 5236 4452 5264
rect 4480 5236 5152 5264
rect 5236 5264 5320 5320
rect 5628 5292 5712 5320
rect 6328 5292 6356 5320
rect 6860 5292 6944 5320
rect 7224 5292 7252 5320
rect 7280 5292 7364 5320
rect 7420 5292 7504 5348
rect 7560 5320 7616 5348
rect 7700 5320 7756 5348
rect 7812 5320 7896 5376
rect 7952 5348 8036 5404
rect 8092 5348 8176 5404
rect 8232 5376 8316 5432
rect 8372 5404 8456 5460
rect 8512 5432 8596 5488
rect 8652 5488 8736 5516
rect 8764 5488 9100 5516
rect 9156 5516 9324 5544
rect 9352 5516 9800 5544
rect 9940 5516 9996 5572
rect 10052 5544 10220 5600
rect 10528 5572 10556 5600
rect 10500 5544 10584 5572
rect 10052 5516 10248 5544
rect 10500 5516 10556 5544
rect 9156 5488 9240 5516
rect 8652 5460 8988 5488
rect 8624 5432 8988 5460
rect 9044 5460 9240 5488
rect 9268 5488 9688 5516
rect 9716 5488 9800 5516
rect 10080 5488 10220 5516
rect 9268 5460 9772 5488
rect 10080 5460 10248 5488
rect 9044 5432 9772 5460
rect 8512 5404 8876 5432
rect 8372 5376 8764 5404
rect 8792 5376 8876 5404
rect 8932 5404 9352 5432
rect 9408 5404 9772 5432
rect 8932 5376 9548 5404
rect 9576 5376 9772 5404
rect 8232 5348 8736 5376
rect 8820 5348 9156 5376
rect 9184 5348 9268 5376
rect 9324 5348 9772 5376
rect 10108 5348 10248 5460
rect 10388 5432 10416 5460
rect 7952 5320 8624 5348
rect 7560 5292 7644 5320
rect 7672 5292 8484 5320
rect 6888 5264 6916 5292
rect 7112 5264 7140 5292
rect 7196 5264 8344 5292
rect 5236 5236 5292 5264
rect 7112 5236 8204 5264
rect 952 5180 1036 5236
rect 2016 5208 2044 5236
rect 3388 5208 3416 5236
rect 4088 5208 4284 5236
rect 4088 5180 4312 5208
rect 4340 5180 4396 5236
rect 4060 5152 4396 5180
rect 4508 5208 4676 5236
rect 4760 5208 5292 5236
rect 7084 5208 7924 5236
rect 4508 5180 4620 5208
rect 4788 5180 5320 5208
rect 5348 5180 5404 5208
rect 4508 5152 4648 5180
rect 1036 5124 1064 5152
rect 4060 5124 4088 5152
rect 4172 5124 4424 5152
rect 4452 5124 4648 5152
rect 4816 5152 4984 5180
rect 5040 5152 5572 5180
rect 6076 5152 6132 5208
rect 6580 5152 6608 5208
rect 6944 5152 7000 5208
rect 7084 5180 7532 5208
rect 7084 5152 7308 5180
rect 4816 5124 4956 5152
rect 1008 5068 1036 5096
rect 1344 5068 1372 5096
rect 1960 5068 2044 5124
rect 3108 5068 3164 5124
rect 3976 5096 4060 5124
rect 3752 5068 3780 5096
rect 3920 5068 4088 5096
rect 4172 5068 4200 5124
rect 616 5012 672 5068
rect 980 5012 1064 5068
rect 1960 5040 2016 5068
rect 2800 5040 2828 5068
rect 3864 5040 4200 5068
rect 4284 5096 4676 5124
rect 4788 5096 4956 5124
rect 2772 5012 2856 5040
rect 3864 5012 4228 5040
rect 4284 5012 4340 5096
rect 4424 5068 4956 5096
rect 5068 5124 5152 5152
rect 5236 5124 5460 5152
rect 5516 5124 5572 5152
rect 7112 5124 7224 5152
rect 7252 5124 7308 5152
rect 7336 5124 7392 5180
rect 7448 5124 7532 5180
rect 7588 5152 7644 5208
rect 7728 5152 7784 5208
rect 7840 5180 7896 5208
rect 7980 5180 8064 5236
rect 8120 5180 8204 5236
rect 8260 5208 8344 5264
rect 8400 5236 8484 5292
rect 8540 5292 8624 5320
rect 8680 5320 8764 5348
rect 8792 5320 9016 5348
rect 8680 5292 9016 5320
rect 9072 5320 9268 5348
rect 9296 5320 9492 5348
rect 9520 5320 9772 5348
rect 9072 5292 9772 5320
rect 10136 5292 10248 5348
rect 8540 5236 8904 5292
rect 8960 5264 9408 5292
rect 9436 5264 9744 5292
rect 8960 5236 9716 5264
rect 10164 5236 10248 5292
rect 10388 5264 10416 5292
rect 8400 5208 8792 5236
rect 8820 5208 9324 5236
rect 9352 5208 9688 5236
rect 8260 5180 8764 5208
rect 8848 5180 9212 5208
rect 9240 5180 9688 5208
rect 10192 5180 10248 5236
rect 7840 5152 7924 5180
rect 7980 5152 8652 5180
rect 7588 5124 7672 5152
rect 7700 5124 8512 5152
rect 5068 5068 5124 5124
rect 5236 5096 5292 5124
rect 952 4900 1120 5012
rect 2800 4984 2828 5012
rect 3892 4984 3920 5012
rect 3948 4984 4340 5012
rect 4452 5040 4984 5068
rect 5040 5040 5124 5068
rect 5236 5040 5264 5068
rect 4452 4984 4480 5040
rect 4508 5012 5180 5040
rect 5208 5012 5292 5040
rect 5376 5012 5432 5124
rect 7112 5096 8372 5124
rect 6104 5068 6132 5096
rect 7084 5068 8008 5096
rect 8148 5068 8232 5096
rect 8288 5068 8344 5096
rect 8428 5068 8512 5124
rect 8568 5124 8652 5152
rect 8708 5152 8792 5180
rect 8820 5152 8932 5180
rect 9016 5152 9212 5180
rect 9268 5152 9436 5180
rect 8708 5124 8848 5152
rect 8876 5124 8932 5152
rect 9100 5124 9212 5152
rect 9240 5124 9436 5152
rect 9492 5124 9716 5180
rect 10164 5152 10248 5180
rect 10192 5124 10248 5152
rect 10360 5124 10388 5152
rect 8568 5096 8820 5124
rect 9100 5096 9352 5124
rect 8540 5068 8792 5096
rect 6132 5040 6188 5068
rect 6804 5040 6888 5068
rect 7084 5040 7812 5068
rect 5544 5012 5600 5040
rect 4508 4984 4620 5012
rect 1764 4928 1792 4984
rect 3780 4956 3808 4984
rect 3864 4956 3892 4984
rect 2212 4928 2240 4956
rect 476 4872 532 4900
rect 476 4844 504 4872
rect 644 4844 700 4900
rect 924 4872 1148 4900
rect 1232 4872 1316 4900
rect 2184 4872 2240 4928
rect 2492 4900 2520 4956
rect 3752 4928 3892 4956
rect 3976 4956 4368 4984
rect 4424 4956 4620 4984
rect 3976 4928 4032 4956
rect 3724 4900 4004 4928
rect 3696 4872 4004 4900
rect 4116 4900 4620 4956
rect 4732 4984 5684 5012
rect 6132 4984 6244 5040
rect 6804 5012 6860 5040
rect 6888 5012 6916 5040
rect 7084 5012 7392 5040
rect 7448 5012 7560 5040
rect 7588 5012 7672 5040
rect 7728 5012 7812 5040
rect 7868 5012 8008 5068
rect 8176 5040 8204 5068
rect 8288 5040 8372 5068
rect 8400 5040 8792 5068
rect 9128 5068 9352 5096
rect 9380 5096 9716 5124
rect 10220 5096 10276 5124
rect 9380 5068 9548 5096
rect 9604 5068 9716 5096
rect 9128 5040 9240 5068
rect 8204 5012 8232 5040
rect 8288 5012 8484 5040
rect 8540 5012 8736 5040
rect 9156 5012 9240 5040
rect 9324 5040 9688 5068
rect 9324 5012 9464 5040
rect 9520 5012 9688 5040
rect 10248 5012 10276 5040
rect 6776 4984 6832 5012
rect 6888 4984 6944 5012
rect 7028 4984 7056 5012
rect 4732 4956 4816 4984
rect 4844 4956 5712 4984
rect 6132 4956 6216 4984
rect 6328 4956 6356 4984
rect 6720 4956 7056 4984
rect 7140 4956 7224 5012
rect 7280 4956 7364 5012
rect 7448 4956 7532 5012
rect 7616 4984 7672 5012
rect 7756 4984 8008 5012
rect 8232 4984 8456 5012
rect 8568 4984 8596 5012
rect 9324 4984 9688 5012
rect 7588 4956 7700 4984
rect 7728 4956 8064 4984
rect 8260 4956 8400 4984
rect 9352 4956 9604 4984
rect 9632 4956 9716 4984
rect 9856 4956 9940 4984
rect 4732 4900 4788 4956
rect 4116 4872 4172 4900
rect 868 4844 896 4872
rect 924 4816 1204 4872
rect 1232 4844 1344 4872
rect 3640 4844 3724 4872
rect 3752 4844 4060 4872
rect 4088 4844 4172 4872
rect 1232 4816 1316 4844
rect 3304 4816 3332 4844
rect 3584 4816 3696 4844
rect 3780 4816 4172 4844
rect 4228 4872 4788 4900
rect 4872 4928 5740 4956
rect 6076 4928 6244 4956
rect 6300 4928 6440 4956
rect 6664 4928 7084 4956
rect 7140 4928 7252 4956
rect 7280 4928 7392 4956
rect 7420 4928 8064 4956
rect 9352 4928 9408 4956
rect 9436 4928 9716 4956
rect 9884 4928 9940 4956
rect 10220 4928 10276 5012
rect 4872 4872 4928 4928
rect 4228 4844 4928 4872
rect 5040 4900 5880 4928
rect 6048 4900 6580 4928
rect 6608 4900 8008 4928
rect 9380 4900 9520 4928
rect 5040 4844 5096 4900
rect 5180 4872 5292 4900
rect 5320 4872 5908 4900
rect 6048 4872 6860 4900
rect 6944 4872 7896 4900
rect 7924 4872 8008 4900
rect 8092 4872 8148 4900
rect 8456 4872 8512 4900
rect 9408 4872 9520 4900
rect 9548 4872 9688 4928
rect 5208 4844 5264 4872
rect 4228 4816 4284 4844
rect 896 4788 1288 4816
rect 868 4760 1260 4788
rect 2156 4760 2240 4816
rect 3528 4788 3724 4816
rect 3780 4788 4284 4816
rect 4368 4816 5096 4844
rect 5180 4816 5264 4844
rect 4368 4788 4452 4816
rect 4508 4788 4592 4816
rect 4620 4788 5264 4816
rect 5348 4788 5404 4872
rect 5488 4844 5572 4872
rect 5516 4788 5572 4844
rect 2744 4760 2772 4788
rect 3500 4760 3836 4788
rect 3920 4760 4424 4788
rect 868 4648 1288 4760
rect 2184 4732 2212 4760
rect 3472 4732 3836 4760
rect 3892 4732 3976 4760
rect 2996 4676 3024 4704
rect 3276 4676 3304 4732
rect 3472 4704 3500 4732
rect 3584 4676 3976 4732
rect 4032 4732 4452 4760
rect 4508 4732 4564 4788
rect 4648 4760 5432 4788
rect 5460 4760 5572 4788
rect 5656 4844 5740 4872
rect 5796 4844 5880 4872
rect 6020 4844 6076 4872
rect 6104 4844 6720 4872
rect 5656 4760 5712 4844
rect 5824 4816 5908 4844
rect 5936 4816 6048 4844
rect 5824 4788 6020 4816
rect 5824 4760 6048 4788
rect 6132 4760 6216 4844
rect 6328 4760 6384 4844
rect 6468 4760 6552 4844
rect 6636 4788 6692 4844
rect 6776 4788 6832 4872
rect 6944 4844 7056 4872
rect 7084 4844 7756 4872
rect 7784 4844 7868 4872
rect 7952 4844 8036 4872
rect 8064 4844 8176 4872
rect 8428 4844 8512 4872
rect 6944 4788 7000 4844
rect 7112 4816 7588 4844
rect 7644 4816 7728 4844
rect 6636 4760 6720 4788
rect 6776 4760 7000 4788
rect 7196 4788 7252 4816
rect 7336 4788 7448 4816
rect 7532 4788 7588 4816
rect 7672 4788 7728 4816
rect 7812 4816 7868 4844
rect 7924 4816 8176 4844
rect 8400 4816 8512 4844
rect 9464 4844 9716 4872
rect 9464 4816 9632 4844
rect 9660 4816 9744 4844
rect 7812 4788 8176 4816
rect 8372 4788 8596 4816
rect 9044 4788 9072 4816
rect 9324 4788 9352 4816
rect 9464 4788 9548 4816
rect 9576 4788 9744 4816
rect 4676 4732 4732 4760
rect 4816 4732 6412 4760
rect 6440 4732 7028 4760
rect 7196 4732 7224 4788
rect 7336 4732 7420 4788
rect 7672 4760 8176 4788
rect 8344 4760 8624 4788
rect 9436 4760 9744 4788
rect 9800 4760 9884 4844
rect 10052 4816 10136 4872
rect 10192 4844 10248 4928
rect 10164 4816 10248 4844
rect 10052 4788 10248 4816
rect 10024 4760 10220 4788
rect 7560 4732 7588 4760
rect 7644 4732 8092 4760
rect 8120 4732 8176 4760
rect 8316 4732 8456 4760
rect 8512 4732 8624 4760
rect 8652 4732 8708 4760
rect 9464 4732 9716 4760
rect 10024 4732 10248 4760
rect 4032 4704 4564 4732
rect 4648 4704 4704 4732
rect 4816 4704 4900 4732
rect 4984 4704 7028 4732
rect 7336 4704 7448 4732
rect 7532 4704 8064 4732
rect 4032 4676 4116 4704
rect 4144 4676 4592 4704
rect 4620 4676 4732 4704
rect 4816 4676 4872 4704
rect 3500 4648 3528 4676
rect 3584 4648 3668 4676
rect 3724 4648 4088 4676
rect 4172 4648 4732 4676
rect 4788 4648 4872 4676
rect 4984 4676 5068 4704
rect 5152 4676 7028 4704
rect 4984 4648 5040 4676
rect 5180 4648 5208 4676
rect 700 4620 756 4648
rect 868 4620 1316 4648
rect 728 4592 756 4620
rect 840 4592 1316 4620
rect 1876 4620 1932 4648
rect 1876 4592 1904 4620
rect 2408 4592 2464 4648
rect 3500 4620 3640 4648
rect 3724 4620 4116 4648
rect 4144 4620 4228 4648
rect 868 4564 1372 4592
rect 2688 4564 2772 4620
rect 3472 4564 3780 4620
rect 3836 4592 4228 4620
rect 4284 4620 4900 4648
rect 4956 4620 5040 4648
rect 5152 4620 5208 4648
rect 4284 4592 4368 4620
rect 4424 4592 5068 4620
rect 5124 4592 5208 4620
rect 5320 4648 5404 4676
rect 5460 4648 6888 4676
rect 5320 4592 5376 4648
rect 5488 4592 5544 4648
rect 5628 4620 5740 4648
rect 5768 4620 6440 4648
rect 6468 4620 6580 4648
rect 6636 4620 6720 4648
rect 6804 4620 6860 4648
rect 3864 4564 4368 4592
rect 4452 4564 5376 4592
rect 5460 4564 5544 4592
rect 5656 4564 5712 4620
rect 5824 4592 5880 4620
rect 5964 4592 6048 4620
rect 6132 4592 6216 4620
rect 5824 4564 5852 4592
rect 868 4536 1400 4564
rect 2688 4536 2744 4564
rect 3248 4536 3276 4564
rect 3528 4536 3808 4564
rect 3836 4536 3920 4564
rect 896 4508 1456 4536
rect 3248 4508 3304 4536
rect 3528 4508 3920 4536
rect 3976 4536 4368 4564
rect 4424 4536 4508 4564
rect 3976 4508 4508 4536
rect 4592 4536 5572 4564
rect 5628 4536 5712 4564
rect 5796 4536 5880 4564
rect 5964 4536 6020 4592
rect 6160 4536 6216 4592
rect 6328 4536 6384 4620
rect 6496 4564 6552 4620
rect 6664 4564 6720 4620
rect 6832 4592 6888 4620
rect 6972 4592 7028 4676
rect 7252 4676 7924 4704
rect 7252 4648 7812 4676
rect 7840 4648 7924 4676
rect 8008 4676 8064 4704
rect 8148 4704 8204 4732
rect 8288 4704 8456 4732
rect 8148 4676 8372 4704
rect 8540 4676 8708 4732
rect 8764 4704 8792 4732
rect 9492 4704 9660 4732
rect 8764 4676 8820 4704
rect 9520 4676 9576 4704
rect 9604 4676 9716 4704
rect 9996 4676 10220 4732
rect 8008 4648 8372 4676
rect 8512 4648 8680 4676
rect 9520 4648 9716 4676
rect 7252 4620 7784 4648
rect 7868 4620 7952 4648
rect 7980 4620 8260 4648
rect 8316 4620 8400 4648
rect 8428 4620 8680 4648
rect 7112 4592 7140 4620
rect 7280 4592 7644 4620
rect 6804 4564 6888 4592
rect 6944 4564 7056 4592
rect 7364 4564 7476 4592
rect 6496 4536 6580 4564
rect 6664 4536 7084 4564
rect 7420 4536 7476 4564
rect 7560 4536 7644 4592
rect 7700 4592 7784 4620
rect 7840 4592 8232 4620
rect 8316 4592 8568 4620
rect 7700 4564 8120 4592
rect 7672 4536 8120 4564
rect 4592 4508 4676 4536
rect 4760 4508 4872 4536
rect 4928 4508 5908 4536
rect 5936 4508 6048 4536
rect 6132 4508 6244 4536
rect 6300 4508 6440 4536
rect 6468 4508 7084 4536
rect 7448 4508 7504 4536
rect 7560 4508 7980 4536
rect 700 4452 756 4508
rect 896 4480 1372 4508
rect 1400 4480 1456 4508
rect 896 4452 1456 4480
rect 1652 4452 1736 4508
rect 616 4424 700 4452
rect 644 4396 700 4424
rect 896 4424 1484 4452
rect 1680 4424 1708 4452
rect 2100 4424 2156 4480
rect 3444 4452 3612 4508
rect 3668 4452 4032 4508
rect 4116 4480 4536 4508
rect 4564 4480 4676 4508
rect 4788 4480 4844 4508
rect 4116 4452 4676 4480
rect 4760 4452 4844 4480
rect 2688 4424 2716 4452
rect 3416 4424 3612 4452
rect 3640 4424 3752 4452
rect 3780 4424 4172 4452
rect 896 4396 1456 4424
rect 924 4368 1456 4396
rect 1484 4396 1512 4424
rect 1484 4368 1540 4396
rect 2352 4368 2408 4424
rect 3192 4368 3276 4424
rect 3416 4396 3724 4424
rect 3808 4396 4172 4424
rect 4256 4424 4844 4452
rect 4956 4480 5040 4508
rect 5096 4480 7112 4508
rect 4956 4424 5012 4480
rect 4256 4396 4340 4424
rect 4368 4396 4872 4424
rect 4928 4396 5012 4424
rect 5124 4452 5236 4480
rect 5264 4452 7112 4480
rect 7448 4480 7980 4508
rect 7448 4452 7840 4480
rect 7896 4452 7980 4480
rect 8036 4508 8120 4536
rect 8176 4564 8260 4592
rect 8288 4564 8568 4592
rect 9548 4592 9716 4648
rect 9548 4564 9632 4592
rect 9660 4564 9716 4592
rect 10024 4620 10192 4676
rect 10024 4564 10052 4620
rect 10108 4592 10164 4620
rect 10304 4592 10360 4648
rect 8176 4508 8428 4564
rect 8036 4480 8428 4508
rect 8512 4480 8596 4564
rect 9576 4536 9716 4564
rect 8988 4480 9016 4508
rect 8036 4452 8288 4480
rect 5124 4396 5180 4452
rect 3500 4368 3752 4396
rect 3780 4368 3864 4396
rect 3920 4368 4312 4396
rect 924 4340 1540 4368
rect 3388 4340 3416 4368
rect 3500 4340 3864 4368
rect 3948 4340 4312 4368
rect 4396 4368 5040 4396
rect 5096 4368 5180 4396
rect 5292 4424 5376 4452
rect 5432 4424 6916 4452
rect 7000 4424 7084 4452
rect 5292 4368 5348 4424
rect 5460 4368 5516 4424
rect 4396 4340 4480 4368
rect 924 4284 1120 4340
rect 1148 4284 1540 4340
rect 1848 4284 1876 4340
rect 3388 4312 3444 4340
rect 3472 4312 3556 4340
rect 952 4256 1148 4284
rect 1204 4256 1568 4284
rect 2324 4256 2380 4312
rect 3388 4284 3556 4312
rect 3612 4312 3864 4340
rect 3920 4312 4004 4340
rect 4060 4312 4480 4340
rect 3612 4284 4004 4312
rect 4088 4284 4480 4312
rect 4536 4340 5376 4368
rect 5432 4340 5516 4368
rect 5628 4396 5712 4424
rect 5768 4396 5880 4424
rect 5936 4396 6608 4424
rect 5628 4340 5684 4396
rect 5796 4340 5852 4396
rect 4536 4312 5544 4340
rect 5600 4312 5712 4340
rect 5768 4312 5852 4340
rect 5964 4368 6048 4396
rect 6132 4368 6216 4396
rect 5964 4340 6020 4368
rect 6160 4340 6216 4368
rect 5964 4312 6048 4340
rect 4536 4284 4648 4312
rect 4676 4284 5908 4312
rect 5936 4284 6048 4312
rect 6132 4312 6216 4340
rect 6328 4368 6412 4396
rect 6496 4368 6580 4396
rect 6328 4340 6384 4368
rect 6524 4340 6580 4368
rect 6328 4312 6412 4340
rect 6496 4312 6580 4340
rect 6664 4340 6748 4424
rect 6832 4396 6916 4424
rect 6860 4368 6916 4396
rect 7028 4396 7084 4424
rect 7476 4396 7672 4452
rect 7728 4424 7812 4452
rect 7896 4424 8288 4452
rect 8372 4424 8596 4480
rect 8960 4452 9016 4480
rect 9576 4480 9744 4536
rect 10276 4508 10304 4536
rect 9576 4452 9660 4480
rect 9688 4452 9744 4480
rect 10388 4480 10444 4508
rect 10388 4452 10472 4480
rect 7756 4396 8176 4424
rect 8232 4396 8316 4424
rect 8344 4396 8568 4424
rect 8848 4396 8876 4424
rect 9604 4396 9716 4452
rect 10416 4424 10444 4452
rect 7028 4368 7112 4396
rect 7504 4368 7560 4396
rect 7588 4368 7672 4396
rect 7728 4368 8148 4396
rect 8232 4368 8484 4396
rect 8540 4368 8568 4396
rect 9604 4368 9688 4396
rect 6832 4340 6916 4368
rect 7000 4340 7196 4368
rect 7308 4340 7364 4368
rect 7504 4340 8036 4368
rect 8064 4340 8176 4368
rect 8204 4340 8456 4368
rect 8680 4340 8736 4368
rect 6664 4312 6776 4340
rect 6804 4312 7224 4340
rect 7308 4312 7336 4340
rect 7532 4312 8008 4340
rect 8092 4312 8484 4340
rect 8540 4312 8568 4340
rect 6132 4284 6244 4312
rect 6300 4284 6440 4312
rect 6468 4284 7224 4312
rect 7532 4284 7868 4312
rect 3388 4256 3696 4284
rect 952 4228 1596 4256
rect 3444 4228 3696 4256
rect 3752 4256 4032 4284
rect 4060 4256 4144 4284
rect 4200 4256 4648 4284
rect 4704 4256 4816 4284
rect 4872 4256 7224 4284
rect 7588 4256 7728 4284
rect 7756 4256 7868 4284
rect 7924 4284 8036 4312
rect 8064 4284 8344 4312
rect 7924 4256 8344 4284
rect 3752 4228 4144 4256
rect 4228 4228 4788 4256
rect 4872 4228 5012 4256
rect 5040 4228 7112 4256
rect 7140 4228 7224 4256
rect 7616 4228 7700 4256
rect 952 4200 1624 4228
rect 952 4172 1652 4200
rect 2072 4172 2100 4200
rect 2632 4172 2688 4228
rect 3472 4200 3724 4228
rect 3752 4200 3836 4228
rect 952 4144 1596 4172
rect 1652 4144 1680 4172
rect 2044 4144 2100 4172
rect 2884 4144 2940 4200
rect 3444 4172 3836 4200
rect 980 4116 1708 4144
rect 3388 4116 3528 4172
rect 3584 4144 3836 4172
rect 3892 4200 4172 4228
rect 4200 4200 4284 4228
rect 3892 4172 4284 4200
rect 4368 4200 4816 4228
rect 4872 4200 4984 4228
rect 4368 4172 4452 4200
rect 4508 4172 4984 4200
rect 3892 4144 3976 4172
rect 3584 4116 3976 4144
rect 1008 4088 1708 4116
rect 3164 4088 3220 4116
rect 3388 4088 3556 4116
rect 3584 4088 3668 4116
rect 3724 4088 3976 4116
rect 4032 4116 4452 4172
rect 4536 4144 4648 4172
rect 4676 4144 4984 4172
rect 5068 4144 5152 4228
rect 5236 4200 6944 4228
rect 7000 4200 7084 4228
rect 5264 4172 5320 4200
rect 4536 4116 4620 4144
rect 4032 4088 4116 4116
rect 812 4060 868 4088
rect 532 4032 560 4060
rect 504 3976 560 4032
rect 1008 4004 1736 4088
rect 2324 4032 2352 4060
rect 1036 3976 1736 4004
rect 1820 3976 1876 4032
rect 3136 4004 3248 4088
rect 3416 4060 3668 4088
rect 3752 4060 4116 4088
rect 4200 4088 4620 4116
rect 4704 4116 5152 4144
rect 5236 4116 5320 4172
rect 5432 4172 5516 4200
rect 5600 4172 5712 4200
rect 5768 4172 5880 4200
rect 5908 4172 6608 4200
rect 6664 4172 6776 4200
rect 5432 4116 5488 4172
rect 5600 4144 5684 4172
rect 5600 4116 5656 4144
rect 5796 4116 5852 4172
rect 4704 4088 4788 4116
rect 4844 4088 5348 4116
rect 5404 4088 5516 4116
rect 5600 4088 5684 4116
rect 5768 4088 5852 4116
rect 5964 4144 6048 4172
rect 6132 4144 6244 4172
rect 5964 4088 6020 4144
rect 6160 4088 6216 4144
rect 6328 4088 6412 4172
rect 6524 4088 6580 4172
rect 6692 4116 6776 4172
rect 6860 4116 6944 4200
rect 7028 4172 7084 4200
rect 7168 4172 7224 4228
rect 7336 4172 7364 4228
rect 7644 4200 7700 4228
rect 7784 4228 8204 4256
rect 8260 4228 8344 4256
rect 8400 4284 8484 4312
rect 8512 4284 8568 4312
rect 9576 4284 9604 4340
rect 8400 4256 8456 4284
rect 8512 4256 8540 4284
rect 8400 4228 8428 4256
rect 7784 4200 8176 4228
rect 8288 4200 8400 4228
rect 7644 4172 8064 4200
rect 8120 4172 8204 4200
rect 8260 4172 8372 4200
rect 10192 4172 10248 4200
rect 7028 4144 7112 4172
rect 7168 4144 7252 4172
rect 7672 4144 8036 4172
rect 8120 4144 8344 4172
rect 9660 4144 9716 4172
rect 10220 4144 10248 4172
rect 7000 4116 7280 4144
rect 7672 4116 7896 4144
rect 6692 4088 6804 4116
rect 6832 4088 7308 4116
rect 7700 4088 7756 4116
rect 7812 4088 7896 4116
rect 7980 4116 8064 4144
rect 8120 4116 8316 4144
rect 9632 4116 9744 4144
rect 7980 4088 8288 4116
rect 9604 4088 9744 4116
rect 4200 4060 4284 4088
rect 4340 4060 4648 4088
rect 4676 4060 4788 4088
rect 3444 4032 3668 4060
rect 3724 4032 3808 4060
rect 3864 4032 4144 4060
rect 4172 4032 4256 4060
rect 4368 4032 4788 4060
rect 4872 4060 5712 4088
rect 5740 4060 5880 4088
rect 5936 4060 6048 4088
rect 6132 4060 6244 4088
rect 6328 4060 6440 4088
rect 6496 4060 7308 4088
rect 4872 4032 4956 4060
rect 5040 4032 7308 4060
rect 7840 4060 7896 4088
rect 7952 4060 8232 4088
rect 8876 4060 8904 4088
rect 9632 4060 9716 4088
rect 7840 4032 8204 4060
rect 3444 4004 3780 4032
rect 3864 4004 4284 4032
rect 4340 4004 4424 4032
rect 1036 3948 1428 3976
rect 1456 3948 1736 3976
rect 1848 3948 1876 3976
rect 2576 3948 2660 3976
rect 3444 3948 3500 4004
rect 3556 3976 3808 4004
rect 3864 3976 3948 4004
rect 4032 3976 4424 4004
rect 4508 4004 4984 4032
rect 5040 4004 5152 4032
rect 4508 3976 4620 4004
rect 4676 3976 5152 4004
rect 5208 4004 7140 4032
rect 5208 3976 5320 4004
rect 3556 3948 3920 3976
rect 4032 3948 4116 3976
rect 4144 3948 4452 3976
rect 4508 3948 4592 3976
rect 1064 3920 1344 3948
rect 1372 3920 1596 3948
rect 1652 3920 1736 3948
rect 2576 3920 2632 3948
rect 3444 3920 3640 3948
rect 1064 3864 1512 3920
rect 1540 3892 1596 3920
rect 1624 3892 1736 3920
rect 2856 3892 2884 3920
rect 3416 3892 3640 3920
rect 3696 3920 3948 3948
rect 4004 3920 4088 3948
rect 3696 3892 4088 3920
rect 4172 3920 4592 3948
rect 4676 3948 5320 3976
rect 5376 3976 5516 4004
rect 5376 3948 5488 3976
rect 5544 3948 5684 4004
rect 5712 3976 6972 4004
rect 5712 3948 6776 3976
rect 4676 3920 4760 3948
rect 4844 3920 5824 3948
rect 5936 3920 6048 3948
rect 6132 3920 6244 3948
rect 6300 3920 6412 3948
rect 6496 3920 6608 3948
rect 4172 3892 4256 3920
rect 4312 3892 4788 3920
rect 4844 3892 4956 3920
rect 1540 3864 1736 3892
rect 2044 3864 2072 3892
rect 3444 3864 3668 3892
rect 3696 3864 3780 3892
rect 3836 3864 4116 3892
rect 4144 3864 4228 3892
rect 4340 3864 4424 3892
rect 4452 3864 4956 3892
rect 5012 3892 5824 3920
rect 5012 3864 5124 3892
rect 1092 3836 1428 3864
rect 1456 3836 1736 3864
rect 3472 3836 3780 3864
rect 3864 3836 4256 3864
rect 4340 3836 4396 3864
rect 1092 3808 1596 3836
rect 1652 3808 1764 3836
rect 3556 3808 3780 3836
rect 3836 3808 3920 3836
rect 1120 3780 1624 3808
rect 1652 3780 1792 3808
rect 868 3752 896 3780
rect 952 3752 1008 3780
rect 1120 3752 1512 3780
rect 1540 3752 1708 3780
rect 1736 3752 1820 3780
rect 2268 3752 2352 3780
rect 3108 3752 3164 3808
rect 3556 3780 3920 3808
rect 4004 3808 4396 3836
rect 4508 3836 4956 3864
rect 4984 3836 5124 3864
rect 5208 3864 5824 3892
rect 5964 3864 6020 3920
rect 6160 3864 6216 3920
rect 5208 3836 5292 3864
rect 4508 3808 4564 3836
rect 4004 3780 4424 3808
rect 4480 3780 4564 3808
rect 4676 3808 5292 3836
rect 5376 3836 5824 3864
rect 5936 3836 6020 3864
rect 6132 3836 6216 3864
rect 6328 3892 6412 3920
rect 6328 3864 6384 3892
rect 6524 3864 6580 3920
rect 6692 3892 6776 3948
rect 6860 3920 6944 3976
rect 7028 3948 7112 4004
rect 7196 3976 7280 4032
rect 7812 4004 8092 4032
rect 8148 4004 8204 4032
rect 7756 3976 8064 4004
rect 8260 3976 8344 4060
rect 9352 4004 9464 4032
rect 8596 3976 8624 4004
rect 9324 3976 9492 4004
rect 9800 3976 9828 4004
rect 7196 3948 7308 3976
rect 7700 3948 7952 3976
rect 7980 3948 8064 3976
rect 8288 3948 8316 3976
rect 8428 3948 8456 3976
rect 9324 3948 9464 3976
rect 7028 3920 7140 3948
rect 7168 3920 7392 3948
rect 7700 3920 7924 3948
rect 8008 3920 8120 3948
rect 8428 3920 8484 3948
rect 9352 3920 9464 3948
rect 6860 3892 6972 3920
rect 7000 3892 7392 3920
rect 7728 3892 7784 3920
rect 7812 3892 7896 3920
rect 8008 3892 8092 3920
rect 6692 3864 6804 3892
rect 6832 3864 7392 3892
rect 7840 3864 7924 3892
rect 7980 3864 8064 3892
rect 6328 3836 6412 3864
rect 6496 3836 6608 3864
rect 6664 3836 7420 3864
rect 7840 3836 8008 3864
rect 8288 3836 8344 3920
rect 8428 3892 8456 3920
rect 9240 3864 9324 3920
rect 9380 3892 9436 3920
rect 9772 3892 9884 3976
rect 10108 3920 10136 3948
rect 9772 3864 9856 3892
rect 5376 3808 5488 3836
rect 5544 3808 5684 3836
rect 5712 3808 5852 3836
rect 5908 3808 6048 3836
rect 6104 3808 6244 3836
rect 6300 3808 7308 3836
rect 7392 3808 7448 3836
rect 7840 3808 7980 3836
rect 4676 3780 4760 3808
rect 4844 3780 7140 3808
rect 7196 3780 7280 3808
rect 3528 3752 3612 3780
rect 3668 3752 3920 3780
rect 3976 3752 4060 3780
rect 868 3724 924 3752
rect 1120 3724 1708 3752
rect 1764 3724 1876 3752
rect 1148 3696 1904 3724
rect 2240 3696 2380 3752
rect 2828 3724 2884 3752
rect 3556 3724 3612 3752
rect 3696 3724 4060 3752
rect 4144 3752 4564 3780
rect 4648 3752 4732 3780
rect 4144 3724 4256 3752
rect 4284 3724 4732 3752
rect 4844 3724 4928 3780
rect 3612 3696 3640 3724
rect 3668 3696 3752 3724
rect 3808 3696 4088 3724
rect 4144 3696 4228 3724
rect 1148 3668 1624 3696
rect 1652 3668 1820 3696
rect 1848 3668 1932 3696
rect 2268 3668 2352 3696
rect 3388 3668 3416 3696
rect 3640 3668 3752 3696
rect 3836 3668 4228 3696
rect 4312 3696 4928 3724
rect 5012 3752 6972 3780
rect 7028 3752 7112 3780
rect 5012 3696 5096 3752
rect 5208 3696 5292 3752
rect 5348 3724 6776 3752
rect 6860 3724 6944 3752
rect 4312 3668 4396 3696
rect 1176 3640 1820 3668
rect 1876 3640 1932 3668
rect 2296 3640 2324 3668
rect 1176 3612 1708 3640
rect 1204 3584 1708 3612
rect 1764 3584 1932 3640
rect 3108 3612 3136 3668
rect 3640 3640 3780 3668
rect 3808 3640 3920 3668
rect 3976 3640 4256 3668
rect 4284 3640 4396 3668
rect 3668 3612 3892 3640
rect 3976 3612 4396 3640
rect 4480 3668 4956 3696
rect 4984 3668 5096 3696
rect 5180 3668 5264 3696
rect 5376 3668 5460 3724
rect 4480 3612 4564 3668
rect 4620 3640 5292 3668
rect 5348 3640 5460 3668
rect 5572 3696 5656 3724
rect 5572 3640 5628 3696
rect 1204 3556 1932 3584
rect 1988 3556 2044 3612
rect 2548 3584 2604 3612
rect 3668 3584 3920 3612
rect 3976 3584 4060 3612
rect 4116 3584 4564 3612
rect 4648 3612 5488 3640
rect 5516 3612 5656 3640
rect 5740 3612 5824 3724
rect 5936 3612 6020 3724
rect 6104 3696 6244 3724
rect 6300 3696 6412 3724
rect 6496 3696 6580 3724
rect 6132 3668 6216 3696
rect 6132 3640 6188 3668
rect 6328 3640 6384 3696
rect 6524 3640 6580 3696
rect 6692 3640 6776 3724
rect 6888 3668 6944 3724
rect 7056 3696 7112 3752
rect 7224 3752 7280 3780
rect 7392 3780 7504 3808
rect 7840 3780 7924 3808
rect 10108 3780 10136 3808
rect 7392 3752 7560 3780
rect 7756 3752 7812 3780
rect 10108 3752 10164 3780
rect 7224 3724 7308 3752
rect 7392 3724 7616 3752
rect 8372 3724 8428 3752
rect 7224 3696 7616 3724
rect 7056 3668 7672 3696
rect 8148 3668 8232 3696
rect 6860 3640 7728 3668
rect 8064 3640 8260 3668
rect 8344 3640 8456 3724
rect 8876 3696 8904 3724
rect 6132 3612 6216 3640
rect 6328 3612 6412 3640
rect 6496 3612 6608 3640
rect 6692 3612 7616 3640
rect 7700 3612 7728 3640
rect 8008 3612 8232 3640
rect 8372 3612 8400 3640
rect 9996 3612 10024 3668
rect 4648 3584 4732 3612
rect 3668 3556 4060 3584
rect 4144 3556 4732 3584
rect 4816 3584 6048 3612
rect 6104 3584 6244 3612
rect 6300 3584 6440 3612
rect 6468 3584 7476 3612
rect 7532 3584 7616 3612
rect 7728 3584 7756 3612
rect 7924 3584 8232 3612
rect 4816 3556 4900 3584
rect 1064 3500 1092 3528
rect 1232 3500 1820 3556
rect 1876 3528 1960 3556
rect 3668 3528 3752 3556
rect 1876 3500 1988 3528
rect 3696 3500 3752 3528
rect 3808 3528 4060 3556
rect 4116 3528 4200 3556
rect 3808 3500 4200 3528
rect 4284 3528 4732 3556
rect 4788 3528 4900 3556
rect 4284 3500 4396 3528
rect 4424 3500 4900 3528
rect 4984 3556 5096 3584
rect 5152 3556 7308 3584
rect 4984 3500 5068 3556
rect 1232 3472 1736 3500
rect 1764 3472 2016 3500
rect 1260 3444 1708 3472
rect 1764 3444 1932 3472
rect 1288 3416 1932 3444
rect 1988 3444 2072 3472
rect 2268 3444 2296 3500
rect 2800 3472 2856 3500
rect 3808 3472 3920 3500
rect 3948 3472 4368 3500
rect 3808 3444 3892 3472
rect 3976 3444 4368 3472
rect 4452 3472 5068 3500
rect 5180 3528 5264 3556
rect 5348 3528 7140 3556
rect 7196 3528 7280 3556
rect 5180 3472 5236 3528
rect 4452 3444 4536 3472
rect 1988 3416 2100 3444
rect 3836 3416 3892 3444
rect 3948 3416 4060 3444
rect 4116 3416 4536 3444
rect 4620 3444 5236 3472
rect 5348 3444 5432 3528
rect 4620 3416 4704 3444
rect 1260 3388 2128 3416
rect 3080 3388 3108 3416
rect 3864 3388 4032 3416
rect 4116 3388 4564 3416
rect 4592 3388 4704 3416
rect 1288 3360 1820 3388
rect 1876 3360 2044 3388
rect 1316 3332 2044 3360
rect 2100 3360 2128 3388
rect 3892 3360 4060 3388
rect 2100 3332 2156 3360
rect 4088 3332 4200 3388
rect 4256 3360 4704 3388
rect 4788 3416 5432 3444
rect 5544 3500 5656 3528
rect 5684 3500 6944 3528
rect 7028 3500 7112 3528
rect 5544 3472 5628 3500
rect 5740 3472 5824 3500
rect 5908 3472 6020 3500
rect 6104 3472 6244 3500
rect 6300 3472 6440 3500
rect 6468 3472 6608 3500
rect 6692 3472 6776 3500
rect 5544 3416 5600 3472
rect 5740 3416 5796 3472
rect 5936 3444 6020 3472
rect 6132 3444 6216 3472
rect 4788 3388 4900 3416
rect 4928 3388 5628 3416
rect 5712 3388 5824 3416
rect 5936 3388 5992 3444
rect 6132 3388 6188 3444
rect 6328 3388 6384 3472
rect 6524 3388 6580 3472
rect 6692 3416 6748 3472
rect 6888 3416 6944 3500
rect 7056 3444 7112 3500
rect 7224 3472 7280 3528
rect 7392 3500 7448 3584
rect 7560 3528 7616 3584
rect 7700 3528 7756 3584
rect 7812 3556 8232 3584
rect 7784 3528 8120 3556
rect 7532 3500 8092 3528
rect 8204 3500 8232 3556
rect 9716 3500 9772 3528
rect 7364 3472 7952 3500
rect 8036 3472 8092 3500
rect 7224 3444 7812 3472
rect 7840 3444 7924 3472
rect 8036 3444 8120 3472
rect 8148 3444 8176 3472
rect 8876 3444 8904 3472
rect 9380 3444 9436 3500
rect 9688 3472 9772 3500
rect 9968 3472 9996 3500
rect 7028 3416 7784 3444
rect 6692 3388 6776 3416
rect 6860 3388 7644 3416
rect 7700 3388 7784 3416
rect 4788 3360 4872 3388
rect 4256 3332 4368 3360
rect 4424 3332 4872 3360
rect 4956 3360 5040 3388
rect 5096 3360 5852 3388
rect 5880 3360 6020 3388
rect 6104 3360 6216 3388
rect 6300 3360 6412 3388
rect 6496 3360 6636 3388
rect 6664 3360 7476 3388
rect 7532 3360 7616 3388
rect 7728 3360 7784 3388
rect 7868 3416 7952 3444
rect 8008 3416 8176 3444
rect 9660 3416 9772 3472
rect 7868 3388 8148 3416
rect 8344 3388 8428 3416
rect 7868 3360 8120 3388
rect 4956 3332 5012 3360
rect 5124 3332 5236 3360
rect 5292 3332 7308 3360
rect 7364 3332 7448 3360
rect 1316 3304 1736 3332
rect 1792 3304 1960 3332
rect 1344 3276 1736 3304
rect 1820 3276 1960 3304
rect 1372 3248 1960 3276
rect 1988 3304 2156 3332
rect 2268 3304 2296 3332
rect 3332 3304 3388 3332
rect 4144 3304 4340 3332
rect 4424 3304 4508 3332
rect 4676 3304 5012 3332
rect 1988 3276 2184 3304
rect 4144 3276 4368 3304
rect 4620 3276 4648 3304
rect 4816 3276 5012 3304
rect 5152 3276 5208 3332
rect 5320 3304 5460 3332
rect 5488 3304 7280 3332
rect 1988 3248 2212 3276
rect 2520 3248 2548 3276
rect 3612 3248 3668 3276
rect 1372 3220 2072 3248
rect 1400 3192 1876 3220
rect 1904 3192 2072 3220
rect 2100 3220 2268 3248
rect 2492 3220 2576 3248
rect 3584 3220 3696 3248
rect 4592 3220 4676 3276
rect 4872 3248 5040 3276
rect 5124 3248 5208 3276
rect 5348 3248 5404 3304
rect 5516 3276 5628 3304
rect 5712 3276 6972 3304
rect 4900 3220 5236 3248
rect 5320 3220 5404 3248
rect 5544 3220 5600 3276
rect 5712 3248 5796 3276
rect 5908 3248 6020 3276
rect 6104 3248 6216 3276
rect 6272 3248 6412 3276
rect 6468 3248 6608 3276
rect 6664 3248 6776 3276
rect 2100 3192 2324 3220
rect 2520 3192 2576 3220
rect 2772 3192 2828 3220
rect 1400 3164 2184 3192
rect 1428 3136 1960 3164
rect 2016 3136 2184 3164
rect 2212 3164 2352 3192
rect 2800 3164 2828 3192
rect 3584 3164 3724 3220
rect 4620 3192 4648 3220
rect 4928 3192 5432 3220
rect 5516 3192 5600 3220
rect 5740 3192 5796 3248
rect 5936 3192 5992 3248
rect 6132 3192 6188 3248
rect 6300 3220 6384 3248
rect 6496 3220 6580 3248
rect 4956 3164 5628 3192
rect 5712 3164 5796 3192
rect 5908 3164 5992 3192
rect 6104 3164 6188 3192
rect 6328 3164 6384 3220
rect 6524 3192 6580 3220
rect 6496 3164 6580 3192
rect 6692 3192 6748 3248
rect 6860 3192 6944 3276
rect 7028 3220 7112 3304
rect 7224 3248 7280 3304
rect 7392 3276 7448 3332
rect 7560 3332 7616 3360
rect 7560 3304 7644 3332
rect 7700 3304 8092 3360
rect 8316 3332 8456 3388
rect 8652 3332 8680 3388
rect 9268 3360 9324 3416
rect 9520 3388 9548 3416
rect 9716 3388 9744 3416
rect 8316 3304 8372 3332
rect 8400 3304 8456 3332
rect 9156 3304 9212 3332
rect 7532 3276 8064 3304
rect 8316 3276 8428 3304
rect 9128 3276 9212 3304
rect 9408 3276 9436 3332
rect 7364 3248 7952 3276
rect 8008 3248 8036 3276
rect 8372 3248 8400 3276
rect 9156 3248 9184 3276
rect 7196 3220 7812 3248
rect 7028 3192 7784 3220
rect 6692 3164 6776 3192
rect 6832 3164 7644 3192
rect 7672 3164 7784 3192
rect 7840 3192 7952 3248
rect 8120 3192 8148 3248
rect 9296 3220 9324 3248
rect 8876 3192 8932 3220
rect 7840 3164 7980 3192
rect 2212 3136 2380 3164
rect 3612 3136 3696 3164
rect 3892 3136 3920 3164
rect 5068 3136 5824 3164
rect 5880 3136 6020 3164
rect 6076 3136 6216 3164
rect 6300 3136 6412 3164
rect 6496 3136 6608 3164
rect 6664 3136 7616 3164
rect 7700 3136 7924 3164
rect 1428 3108 1988 3136
rect 2016 3108 2296 3136
rect 2324 3108 2436 3136
rect 3024 3108 3080 3136
rect 5124 3108 5208 3136
rect 5292 3108 7448 3136
rect 1456 3080 2100 3108
rect 1316 3024 1344 3052
rect 1484 3024 1904 3080
rect 1932 3052 2072 3080
rect 2128 3052 2296 3108
rect 2352 3080 2464 3108
rect 3052 3080 3080 3108
rect 4144 3080 4172 3108
rect 2324 3052 2520 3080
rect 2772 3052 2828 3080
rect 1932 3024 2408 3052
rect 1512 2996 2016 3024
rect 1540 2968 2016 2996
rect 2044 2996 2184 3024
rect 2240 2996 2408 3024
rect 2464 3024 2576 3052
rect 2772 3024 2856 3052
rect 3612 3024 3640 3052
rect 4648 3024 4676 3052
rect 5124 3024 5180 3108
rect 5320 3080 5404 3108
rect 5488 3080 7280 3108
rect 2464 2996 2632 3024
rect 2800 2996 2828 3024
rect 3276 2996 3332 3024
rect 4620 2996 4704 3024
rect 5124 2996 5208 3024
rect 5320 2996 5376 3080
rect 5516 3052 5600 3080
rect 5684 3052 6972 3080
rect 7000 3052 7112 3080
rect 2044 2968 2212 2996
rect 2240 2968 2520 2996
rect 1540 2940 2296 2968
rect 1568 2912 1932 2940
rect 1960 2912 2100 2940
rect 2156 2912 2296 2940
rect 2352 2940 2520 2968
rect 2576 2940 2632 2996
rect 2352 2912 2632 2940
rect 3024 2912 3080 2968
rect 1568 2884 2436 2912
rect 1596 2856 2212 2884
rect 2268 2856 2436 2884
rect 2464 2884 2632 2912
rect 3248 2884 3360 2996
rect 4620 2968 4732 2996
rect 4984 2968 5012 2996
rect 5096 2968 5236 2996
rect 5264 2968 5404 2996
rect 5516 2968 5572 3052
rect 5712 3024 5796 3052
rect 5908 3024 5992 3052
rect 6076 3024 6216 3052
rect 6272 3024 6412 3052
rect 6468 3024 6608 3052
rect 6664 3024 6776 3052
rect 6832 3024 6944 3052
rect 5712 2968 5768 3024
rect 4620 2940 4704 2968
rect 4956 2912 5040 2968
rect 5068 2940 5600 2968
rect 5684 2940 5796 2968
rect 5908 2940 5964 3024
rect 6104 2996 6188 3024
rect 6300 2996 6384 3024
rect 6496 2996 6580 3024
rect 6104 2968 6160 2996
rect 6300 2968 6356 2996
rect 6496 2968 6552 2996
rect 6692 2968 6748 3024
rect 6860 2968 6944 3024
rect 7028 2996 7112 3052
rect 7196 3052 7280 3080
rect 7364 3080 7448 3108
rect 7532 3108 7616 3136
rect 7672 3108 7896 3136
rect 8904 3108 8988 3136
rect 9184 3108 9212 3164
rect 9772 3136 9800 3164
rect 9436 3108 9464 3136
rect 7532 3080 7868 3108
rect 8876 3080 8988 3108
rect 7364 3052 7784 3080
rect 8652 3052 8736 3080
rect 8904 3052 8988 3080
rect 9296 3052 9352 3108
rect 9408 3080 9492 3108
rect 9408 3052 9464 3080
rect 7196 3024 7308 3052
rect 7336 3024 7784 3052
rect 8624 3024 8764 3052
rect 8904 3024 8960 3052
rect 9296 3024 9324 3052
rect 7168 2996 7644 3024
rect 7672 2996 7784 3024
rect 8400 2996 8428 3024
rect 7000 2968 7616 2996
rect 6104 2940 6188 2968
rect 6300 2940 6384 2968
rect 6496 2940 6580 2968
rect 6664 2940 6776 2968
rect 6832 2940 7448 2968
rect 5068 2912 5824 2940
rect 5880 2912 5992 2940
rect 6076 2912 6188 2940
rect 6272 2912 6384 2940
rect 6468 2912 7280 2940
rect 2464 2856 2660 2884
rect 3612 2856 3640 2912
rect 5096 2856 5180 2912
rect 5264 2884 7112 2912
rect 1624 2828 2716 2856
rect 5124 2828 5180 2856
rect 5292 2856 5404 2884
rect 5460 2856 6944 2884
rect 5292 2828 5376 2856
rect 5488 2828 5600 2856
rect 5684 2828 5824 2856
rect 5852 2828 6580 2856
rect 6608 2828 6748 2856
rect 1624 2800 2128 2828
rect 1456 2772 1484 2800
rect 1652 2772 2128 2800
rect 2184 2800 2352 2828
rect 2380 2800 2548 2828
rect 2604 2800 2772 2828
rect 3864 2800 3892 2828
rect 5180 2800 5404 2828
rect 5488 2800 5572 2828
rect 5684 2800 5796 2828
rect 2184 2772 2800 2800
rect 3612 2772 3668 2800
rect 5180 2772 5600 2800
rect 5656 2772 5796 2800
rect 5880 2772 5992 2828
rect 1680 2744 2464 2772
rect 1680 2716 2268 2744
rect 2296 2716 2464 2744
rect 2492 2716 2744 2772
rect 2772 2716 2828 2772
rect 1512 2688 1540 2716
rect 1708 2688 2352 2716
rect 2380 2688 2576 2716
rect 1736 2660 2380 2688
rect 2408 2660 2576 2688
rect 2604 2688 2828 2716
rect 2604 2660 2744 2688
rect 3164 2660 3248 2744
rect 3584 2716 3696 2772
rect 4900 2744 4928 2772
rect 5180 2744 5824 2772
rect 5852 2744 5992 2772
rect 6076 2744 6188 2828
rect 6272 2772 6384 2828
rect 6440 2800 6552 2828
rect 6468 2772 6552 2800
rect 6636 2800 6748 2828
rect 6832 2828 6916 2856
rect 7000 2828 7112 2884
rect 7168 2884 7280 2912
rect 7336 2912 7448 2940
rect 7504 2940 7616 2968
rect 7672 2968 7756 2996
rect 7672 2940 7728 2968
rect 8064 2940 8148 2996
rect 8596 2968 8764 3024
rect 8624 2940 8764 2968
rect 9184 2940 9212 2996
rect 7504 2912 7700 2940
rect 8092 2912 8120 2940
rect 8624 2912 8736 2940
rect 7336 2884 7672 2912
rect 8848 2884 8876 2940
rect 9100 2912 9128 2940
rect 7168 2856 7644 2884
rect 9072 2856 9128 2912
rect 7140 2828 7616 2856
rect 6832 2800 6944 2828
rect 6972 2800 7448 2828
rect 7476 2800 7532 2828
rect 6636 2772 7280 2800
rect 7308 2772 7420 2800
rect 8344 2772 8400 2828
rect 6244 2744 6384 2772
rect 6440 2744 7252 2772
rect 7336 2744 7448 2772
rect 9100 2744 9156 2772
rect 4900 2716 4956 2744
rect 5180 2716 5208 2744
rect 5236 2716 6916 2744
rect 3612 2688 3668 2716
rect 5264 2688 5404 2716
rect 5460 2688 6748 2716
rect 6776 2688 6916 2716
rect 1736 2632 2296 2660
rect 2324 2632 2716 2660
rect 3836 2632 3892 2688
rect 5264 2660 5376 2688
rect 5460 2660 5572 2688
rect 4648 2632 4676 2660
rect 5180 2632 5208 2660
rect 5264 2632 5404 2660
rect 5432 2632 5572 2660
rect 5656 2660 5796 2688
rect 5852 2660 6020 2688
rect 6048 2660 6384 2688
rect 6412 2660 6552 2688
rect 5656 2632 5768 2660
rect 5880 2632 5992 2660
rect 1764 2604 2492 2632
rect 2520 2604 2716 2632
rect 4116 2604 4144 2632
rect 5180 2604 5236 2632
rect 5264 2604 5796 2632
rect 5852 2604 5992 2632
rect 6048 2632 6160 2660
rect 6048 2604 6188 2632
rect 6244 2604 6356 2660
rect 6440 2632 6552 2660
rect 6608 2660 6720 2688
rect 6804 2660 6916 2688
rect 6972 2688 7084 2744
rect 7168 2716 7448 2744
rect 7140 2688 7420 2716
rect 9072 2688 9184 2744
rect 9464 2716 9492 2744
rect 6972 2660 7392 2688
rect 9072 2660 9156 2688
rect 6608 2632 6748 2660
rect 6776 2632 7420 2660
rect 6412 2604 7252 2632
rect 7308 2604 7420 2632
rect 7784 2604 7840 2632
rect 8792 2604 8848 2632
rect 1792 2576 2688 2604
rect 3612 2576 3640 2604
rect 4088 2576 4172 2604
rect 5320 2576 7084 2604
rect 7140 2576 7420 2604
rect 8764 2576 8848 2604
rect 9016 2576 9128 2604
rect 1792 2548 2408 2576
rect 2436 2548 2604 2576
rect 2632 2548 2660 2576
rect 4116 2548 4144 2576
rect 5376 2548 5404 2576
rect 5460 2548 6888 2576
rect 6972 2548 7084 2576
rect 7112 2548 7392 2576
rect 8792 2548 8848 2576
rect 8988 2548 9156 2576
rect 1652 2520 1680 2548
rect 1848 2520 2660 2548
rect 1848 2492 2520 2520
rect 2548 2492 2660 2520
rect 1876 2464 2688 2492
rect 3024 2464 3080 2520
rect 5488 2492 5572 2548
rect 5628 2520 5796 2548
rect 5824 2520 6552 2548
rect 6580 2520 6720 2548
rect 6776 2520 6916 2548
rect 6944 2520 7392 2548
rect 8876 2520 8904 2548
rect 8960 2520 9184 2548
rect 5656 2492 5768 2520
rect 5852 2492 5964 2520
rect 1708 2436 1736 2464
rect 1904 2436 2632 2464
rect 1932 2408 2632 2436
rect 2660 2408 2688 2464
rect 3192 2436 3220 2464
rect 4900 2436 4956 2492
rect 5460 2464 5768 2492
rect 5824 2464 5964 2492
rect 6048 2464 6160 2520
rect 6244 2492 6356 2520
rect 6216 2464 6356 2492
rect 6412 2492 6524 2520
rect 6608 2492 6748 2520
rect 6776 2492 7252 2520
rect 7280 2492 7336 2520
rect 7504 2492 7588 2520
rect 8960 2492 9016 2520
rect 9044 2492 9156 2520
rect 6412 2464 7252 2492
rect 5432 2436 7056 2464
rect 7140 2436 7252 2464
rect 7476 2464 7616 2492
rect 7476 2436 7644 2464
rect 8988 2436 9128 2492
rect 9296 2436 9324 2464
rect 3164 2408 3248 2436
rect 4592 2408 4676 2436
rect 5404 2408 6720 2436
rect 6748 2408 6888 2436
rect 1960 2380 2688 2408
rect 1988 2352 2688 2380
rect 3136 2352 3276 2408
rect 4564 2380 4704 2408
rect 5404 2380 5572 2408
rect 5628 2380 6524 2408
rect 1988 2324 2660 2352
rect 3052 2324 3080 2352
rect 3164 2324 3248 2352
rect 2016 2296 2632 2324
rect 4536 2296 4704 2380
rect 5460 2352 5544 2380
rect 5628 2352 5740 2380
rect 5824 2352 5964 2380
rect 5460 2324 5768 2352
rect 5824 2324 5936 2352
rect 6020 2324 6132 2380
rect 6216 2324 6328 2380
rect 6412 2352 6524 2380
rect 6580 2380 6692 2408
rect 6776 2380 6888 2408
rect 6944 2380 7308 2436
rect 7476 2380 7616 2436
rect 9016 2408 9044 2436
rect 9072 2408 9100 2436
rect 6580 2352 6720 2380
rect 6748 2352 7252 2380
rect 7280 2352 7336 2380
rect 7504 2352 7588 2380
rect 7896 2352 7952 2380
rect 6384 2324 7084 2352
rect 7112 2324 7224 2352
rect 7280 2324 7364 2352
rect 5432 2296 7056 2324
rect 7112 2296 7392 2324
rect 7868 2296 7980 2352
rect 8344 2324 8372 2352
rect 8288 2296 8400 2324
rect 2072 2268 2604 2296
rect 2856 2268 2884 2296
rect 4116 2268 4144 2296
rect 4564 2268 4676 2296
rect 5432 2268 6860 2296
rect 6944 2268 7392 2296
rect 1876 2240 1904 2268
rect 2072 2240 2548 2268
rect 5460 2240 5572 2268
rect 5600 2240 6524 2268
rect 6552 2240 6692 2268
rect 6748 2240 6888 2268
rect 6916 2240 7392 2268
rect 7840 2240 7952 2296
rect 8288 2240 8428 2296
rect 9044 2240 9072 2268
rect 2100 2212 2436 2240
rect 2464 2212 2492 2240
rect 4312 2212 4424 2240
rect 5460 2212 5544 2240
rect 5628 2212 5740 2240
rect 2128 2184 2464 2212
rect 3052 2184 3080 2212
rect 4284 2184 4452 2212
rect 5124 2184 5208 2212
rect 5432 2184 5572 2212
rect 5600 2184 5740 2212
rect 5796 2184 5936 2240
rect 5992 2184 6132 2240
rect 6188 2184 6328 2240
rect 6384 2212 6496 2240
rect 6580 2212 6720 2240
rect 6748 2212 7224 2240
rect 7280 2212 7364 2240
rect 7784 2212 7952 2240
rect 8092 2212 8120 2240
rect 8288 2212 8400 2240
rect 6384 2184 7056 2212
rect 7084 2184 7224 2212
rect 7252 2184 7392 2212
rect 7756 2184 7924 2212
rect 8064 2184 8148 2212
rect 8316 2184 8344 2212
rect 1960 2100 2016 2184
rect 2156 2156 2464 2184
rect 3444 2156 3472 2184
rect 2184 2128 2520 2156
rect 4116 2128 4144 2156
rect 4284 2128 4340 2184
rect 4396 2128 4452 2184
rect 4620 2156 4648 2184
rect 4872 2128 4928 2184
rect 5124 2156 5236 2184
rect 5404 2156 7028 2184
rect 7084 2156 7392 2184
rect 7700 2156 7924 2184
rect 8036 2156 8148 2184
rect 5124 2128 5208 2156
rect 5404 2128 6692 2156
rect 6720 2128 6860 2156
rect 6916 2128 7364 2156
rect 7644 2128 7784 2156
rect 7812 2128 7896 2156
rect 8064 2128 8148 2156
rect 8456 2128 8484 2156
rect 2212 2100 2520 2128
rect 2744 2100 2772 2128
rect 3248 2100 3276 2128
rect 3640 2100 3696 2128
rect 4284 2100 4452 2128
rect 2240 2072 2520 2100
rect 4312 2072 4424 2100
rect 5432 2072 5544 2128
rect 5600 2100 6496 2128
rect 5600 2072 5740 2100
rect 2296 2044 2520 2072
rect 5376 2044 5544 2072
rect 5572 2044 5740 2072
rect 5796 2044 5936 2100
rect 5992 2044 6104 2100
rect 6160 2044 6300 2100
rect 6356 2072 6496 2100
rect 6552 2100 6664 2128
rect 6748 2100 7336 2128
rect 7532 2100 7560 2128
rect 7616 2100 7896 2128
rect 8176 2100 8204 2128
rect 8932 2100 9016 2128
rect 6552 2072 7224 2100
rect 7616 2072 7868 2100
rect 8960 2072 9016 2100
rect 6356 2044 7028 2072
rect 7084 2044 7196 2072
rect 2324 2016 2520 2044
rect 3472 2016 3500 2044
rect 4620 2016 4648 2044
rect 5376 2016 6832 2044
rect 2352 1988 2492 2016
rect 3276 1988 3304 2016
rect 2380 1960 2548 1988
rect 3668 1960 3696 1988
rect 4116 1960 4144 2016
rect 4872 1988 4928 2016
rect 5152 1960 5180 2016
rect 5404 1988 6664 2016
rect 5404 1960 5544 1988
rect 5572 1960 6300 1988
rect 6328 1960 6468 1988
rect 2184 1932 2212 1960
rect 2408 1932 2548 1960
rect 2436 1904 2576 1932
rect 3892 1904 3920 1932
rect 4368 1904 4396 1960
rect 5292 1932 5516 1960
rect 5600 1932 5712 1960
rect 5796 1932 5908 1960
rect 5292 1904 5740 1932
rect 5768 1904 5908 1932
rect 5964 1904 6104 1960
rect 6160 1932 6272 1960
rect 6356 1932 6468 1960
rect 6524 1960 6664 1988
rect 6720 1988 6832 2016
rect 6888 2016 7196 2044
rect 7616 2016 7756 2072
rect 7784 2016 7840 2072
rect 6888 1988 7168 2016
rect 6720 1960 7168 1988
rect 7532 1988 7840 2016
rect 7532 1960 7700 1988
rect 7728 1960 7812 1988
rect 6524 1932 7056 1960
rect 7588 1932 7700 1960
rect 7756 1932 7784 1960
rect 6160 1904 7000 1932
rect 7448 1904 7532 1932
rect 7588 1904 7784 1932
rect 8512 1904 8540 1932
rect 8792 1904 8820 1932
rect 2464 1876 2604 1904
rect 3500 1876 3528 1904
rect 4620 1876 4648 1904
rect 5292 1876 6832 1904
rect 6860 1876 6972 1904
rect 7420 1876 7784 1904
rect 8764 1876 8820 1904
rect 2492 1848 2604 1876
rect 4144 1848 4172 1876
rect 4872 1848 4900 1876
rect 2520 1820 2660 1848
rect 5152 1820 5180 1876
rect 5404 1848 6468 1876
rect 6496 1848 6636 1876
rect 6692 1848 6972 1876
rect 7448 1848 7644 1876
rect 7672 1848 7756 1876
rect 8204 1848 8232 1876
rect 5404 1820 5516 1848
rect 2548 1764 2576 1820
rect 2632 1792 2688 1820
rect 4368 1792 4424 1820
rect 5348 1792 5516 1820
rect 5572 1792 5712 1848
rect 5768 1820 6104 1848
rect 5768 1792 5908 1820
rect 5964 1792 6076 1820
rect 6132 1792 6272 1848
rect 6328 1820 6440 1848
rect 6496 1820 6972 1848
rect 7420 1820 7700 1848
rect 6328 1792 6804 1820
rect 6832 1792 6944 1820
rect 7420 1792 7644 1820
rect 7952 1792 7980 1820
rect 2660 1764 2688 1792
rect 3360 1764 3388 1792
rect 3920 1764 3948 1792
rect 4620 1764 4648 1792
rect 5348 1764 6636 1792
rect 4872 1736 4928 1764
rect 5488 1736 6440 1764
rect 2688 1708 2716 1736
rect 3752 1708 3780 1736
rect 5152 1708 5180 1736
rect 3556 1680 3584 1708
rect 4396 1680 4424 1708
rect 5572 1680 5712 1736
rect 5740 1680 5908 1736
rect 5936 1708 6104 1736
rect 6132 1708 6272 1736
rect 6300 1708 6440 1736
rect 6468 1736 6636 1764
rect 6664 1764 6804 1792
rect 6860 1764 6944 1792
rect 7448 1764 7532 1792
rect 6664 1736 6916 1764
rect 7448 1736 7504 1764
rect 6468 1708 6888 1736
rect 5936 1680 6076 1708
rect 6132 1680 6832 1708
rect 3948 1652 3976 1680
rect 5376 1652 5404 1680
rect 5516 1652 6608 1680
rect 6636 1652 6776 1680
rect 4620 1624 4648 1652
rect 4872 1624 4928 1652
rect 5516 1624 6412 1652
rect 6468 1624 6748 1652
rect 4536 1596 4676 1624
rect 5124 1596 5180 1624
rect 5572 1596 5712 1624
rect 5740 1596 5880 1624
rect 5936 1596 6076 1624
rect 6104 1596 6244 1624
rect 6300 1596 6720 1624
rect 7000 1596 7056 1624
rect 2660 1568 2688 1596
rect 4396 1568 4424 1596
rect 4508 1568 4704 1596
rect 5544 1568 6580 1596
rect 4480 1540 4564 1568
rect 4648 1540 4732 1568
rect 5376 1540 5404 1568
rect 5544 1540 6412 1568
rect 2828 1456 2856 1484
rect 3976 1456 4004 1484
rect 4480 1456 4536 1540
rect 4676 1456 4732 1540
rect 5544 1512 5684 1540
rect 5740 1512 5880 1540
rect 5908 1512 6048 1540
rect 6076 1512 6244 1540
rect 6272 1512 6412 1540
rect 6440 1540 6580 1568
rect 6608 1540 6692 1596
rect 6944 1568 7056 1596
rect 7476 1568 7504 1596
rect 6944 1540 7084 1568
rect 8344 1540 8372 1596
rect 6440 1512 6664 1540
rect 6944 1512 7056 1540
rect 5348 1484 5404 1512
rect 5572 1484 6552 1512
rect 6972 1484 7028 1512
rect 7924 1484 8008 1512
rect 4480 1428 4564 1456
rect 4648 1428 4732 1456
rect 4900 1428 4928 1456
rect 2912 1400 2940 1428
rect 4508 1400 4704 1428
rect 5320 1400 5432 1484
rect 5600 1456 5880 1484
rect 5908 1456 6524 1484
rect 5600 1428 5628 1456
rect 5656 1428 6216 1456
rect 6244 1428 6524 1456
rect 5600 1400 6468 1428
rect 7896 1400 8036 1484
rect 8204 1456 8232 1484
rect 4536 1372 4676 1400
rect 5740 1372 6020 1400
rect 6076 1372 6384 1400
rect 6888 1372 6916 1400
rect 7924 1372 8008 1400
rect 3024 1344 3052 1372
rect 5320 1344 5348 1372
rect 5768 1344 6020 1372
rect 6048 1344 6188 1372
rect 6216 1344 6356 1372
rect 7980 1344 8008 1372
rect 3388 1316 3416 1344
rect 5292 1288 5376 1344
rect 5768 1288 5852 1344
rect 5880 1288 6160 1344
rect 6244 1316 6272 1344
rect 5796 1260 5992 1288
rect 6076 1260 6132 1288
rect 3220 1232 3248 1260
rect 7560 1148 7588 1176
rect 7448 1092 7476 1120
rect 7336 1036 7364 1064
rect 3808 980 3836 1036
rect 5544 980 5628 1008
rect 2828 896 2856 952
rect 5516 924 5628 980
rect 6580 952 6608 980
rect 5544 896 5600 924
rect 4788 868 4816 896
rect 6636 840 6664 868
rect 4704 756 4732 784
rect 4816 728 4844 756
<< end >>
