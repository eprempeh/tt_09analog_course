magic
tech sky130A
timestamp 1771423184
<< metal1 >>
rect 2655 3960 2700 4005
rect 2745 3915 2925 3960
rect 2790 3870 3060 3915
rect 2880 3825 3150 3870
rect 1620 3780 1665 3825
rect 2970 3780 3240 3825
rect 1215 3735 1260 3780
rect 1350 3736 1395 3780
rect 1440 3736 1530 3780
rect 1350 3735 1530 3736
rect 1710 3735 1890 3780
rect 3015 3735 3285 3780
rect 1080 3691 1485 3735
rect 1080 3690 1350 3691
rect 990 3645 1125 3690
rect 1215 3645 1305 3690
rect 1395 3645 1485 3691
rect 1710 3645 2025 3735
rect 3015 3690 3375 3735
rect 3015 3645 3420 3690
rect 900 3600 1035 3645
rect 1350 3600 1440 3645
rect 1620 3600 2070 3645
rect 3060 3600 3465 3645
rect 900 3555 945 3600
rect 1305 3555 1395 3600
rect 1575 3555 2025 3600
rect 3015 3555 3510 3600
rect 855 3510 945 3555
rect 1215 3510 1395 3555
rect 1530 3510 1980 3555
rect 2295 3510 2385 3555
rect 2790 3510 2835 3555
rect 810 3465 900 3510
rect 1080 3465 1125 3510
rect 1215 3465 1260 3510
rect 1440 3465 1935 3510
rect 765 3420 855 3465
rect 1035 3420 1170 3465
rect 720 3375 855 3420
rect 945 3375 1170 3420
rect 1395 3420 1845 3465
rect 2745 3420 2835 3510
rect 3015 3510 3555 3555
rect 3015 3465 3600 3510
rect 2925 3420 3645 3465
rect 1395 3375 1755 3420
rect 2970 3375 3690 3420
rect 675 3330 810 3375
rect 900 3330 1080 3375
rect 630 3285 810 3330
rect 855 3285 1080 3330
rect 1350 3330 1530 3375
rect 2925 3330 3735 3375
rect 1350 3285 1440 3330
rect 2475 3285 2520 3330
rect 2835 3285 3780 3330
rect 630 3240 1080 3285
rect 1755 3240 1800 3285
rect 2385 3240 2655 3285
rect 2790 3240 3825 3285
rect 585 3195 1035 3240
rect 1755 3195 1845 3240
rect 2340 3195 2700 3240
rect 2745 3195 3825 3240
rect 540 3105 1035 3195
rect 2340 3150 2610 3195
rect 2745 3150 3870 3195
rect 2295 3105 2430 3150
rect 2520 3105 2655 3150
rect 2700 3105 3870 3150
rect 495 3060 990 3105
rect 2250 3060 2385 3105
rect 2475 3060 3915 3105
rect 495 3015 810 3060
rect 450 2970 810 3015
rect 450 2925 720 2970
rect 450 2880 675 2925
rect 765 2880 810 2970
rect 900 2925 945 3015
rect 2160 2970 2340 3060
rect 2475 3015 3960 3060
rect 2475 2970 2520 3015
rect 2160 2925 2205 2970
rect 2250 2925 2340 2970
rect 2565 2925 3960 3015
rect 1935 2880 1980 2925
rect 2295 2880 2340 2925
rect 2520 2880 4005 2925
rect 405 2835 585 2880
rect 2475 2835 4005 2880
rect 450 2790 585 2835
rect 1845 2790 1890 2835
rect 450 2745 540 2790
rect 450 2655 495 2745
rect 1935 2700 1980 2790
rect 2475 2745 4050 2835
rect 2115 2700 4050 2745
rect 2070 2655 4050 2700
rect 2025 2610 2295 2655
rect 2340 2610 4095 2655
rect 1935 2565 2160 2610
rect 2205 2565 3105 2610
rect 360 2520 405 2565
rect 1080 2520 1125 2565
rect 1935 2520 3060 2565
rect 3240 2520 4095 2610
rect 315 2475 405 2520
rect 1935 2475 2385 2520
rect 2430 2475 2655 2520
rect 2835 2475 3060 2520
rect 3195 2475 4095 2520
rect 360 2340 405 2475
rect 1755 2430 1845 2475
rect 1890 2431 2250 2475
rect 1890 2430 2115 2431
rect 2160 2430 2250 2431
rect 2295 2430 2610 2475
rect 1755 2385 1980 2430
rect 2205 2385 2250 2430
rect 2340 2385 2610 2430
rect 1710 2340 1935 2385
rect 2430 2340 2610 2385
rect 2925 2430 3060 2475
rect 3240 2430 4050 2475
rect 2925 2385 3105 2430
rect 3285 2385 4050 2430
rect 2925 2340 3150 2385
rect 1710 2295 1890 2340
rect 2295 2295 2340 2340
rect 2430 2295 2520 2340
rect 2700 2295 3150 2340
rect 2430 2250 2475 2295
rect 2610 2250 3150 2295
rect 3285 2295 4095 2385
rect 3285 2250 3960 2295
rect 360 2205 405 2250
rect 2610 2205 3960 2250
rect 4050 2250 4095 2295
rect 1755 2160 2160 2205
rect 1710 2115 2160 2160
rect 2880 2115 3915 2205
rect 4050 2115 4140 2250
rect 1665 2112 2160 2115
rect 1665 2070 2164 2112
rect 1575 2025 2164 2070
rect 2835 2070 3915 2115
rect 4095 2070 4140 2115
rect 2835 2025 3555 2070
rect 3645 2025 3915 2070
rect 360 1980 450 2025
rect 1575 1980 2295 2025
rect 2475 1980 2520 2025
rect 2700 1980 3240 2025
rect 3330 1980 3375 2025
rect 3735 1980 3915 2025
rect 360 1845 540 1980
rect 1485 1935 2385 1980
rect 2430 1935 3285 1980
rect 3780 1935 3915 1980
rect 4050 1935 4095 1980
rect 1440 1890 2790 1935
rect 2925 1890 3015 1935
rect 3060 1890 3285 1935
rect 3330 1890 3465 1935
rect 360 1755 585 1845
rect 1395 1755 2835 1890
rect 2925 1845 3465 1890
rect 2970 1800 3465 1845
rect 3825 1800 3915 1935
rect 4005 1845 4095 1935
rect 3015 1755 3465 1800
rect 3870 1755 3915 1800
rect 360 1710 630 1755
rect 1395 1710 2880 1755
rect 3015 1710 3420 1755
rect 360 1665 675 1710
rect 1395 1665 2925 1710
rect 3060 1665 3375 1710
rect 405 1575 675 1665
rect 1350 1620 2925 1665
rect 1395 1575 2925 1620
rect 3105 1620 3330 1665
rect 3870 1620 3915 1665
rect 3105 1575 3240 1620
rect 405 1530 720 1575
rect 1395 1530 2970 1575
rect 3150 1530 3195 1575
rect 450 1485 720 1530
rect 900 1485 945 1530
rect 1440 1485 3060 1530
rect 450 1440 765 1485
rect 1485 1440 3060 1485
rect 3240 1440 3285 1485
rect 495 1395 810 1440
rect 1485 1395 3285 1440
rect 495 1350 855 1395
rect 1575 1350 3285 1395
rect 540 1305 855 1350
rect 1665 1305 1755 1350
rect 1845 1305 1890 1350
rect 1935 1305 2025 1350
rect 2070 1305 3240 1350
rect 3330 1305 3375 1350
rect 540 1260 945 1305
rect 1440 1260 1485 1305
rect 1980 1260 3195 1305
rect 585 1215 990 1260
rect 2115 1215 3150 1260
rect 630 1170 1035 1215
rect 1305 1170 1350 1215
rect 2025 1170 3105 1215
rect 3465 1170 3510 1215
rect 630 1125 1080 1170
rect 2070 1125 3060 1170
rect 675 1080 1125 1125
rect 2070 1080 3015 1125
rect 720 990 1080 1080
rect 2115 1035 2970 1080
rect 3645 1035 3690 1080
rect 2205 990 2970 1035
rect 3600 990 3690 1035
rect 765 945 1080 990
rect 1260 945 1305 990
rect 810 900 1035 945
rect 1845 900 1890 990
rect 2160 945 2925 990
rect 3015 945 3060 990
rect 2205 900 2970 945
rect 3150 900 3195 945
rect 3330 900 3375 945
rect 855 855 990 900
rect 1755 855 1800 900
rect 2160 855 2970 900
rect 3105 855 3195 900
rect 900 810 1035 855
rect 945 765 1035 810
rect 990 720 1035 765
rect 2160 810 2925 855
rect 3060 810 3150 855
rect 2160 765 2880 810
rect 3015 765 3150 810
rect 2160 720 2790 765
rect 2970 720 3105 765
rect 2205 675 2790 720
rect 2205 630 2700 675
rect 1800 585 1845 630
rect 2250 585 2655 630
rect 2790 585 2835 630
rect 1800 540 1890 585
rect 2295 540 2610 585
rect 2340 495 2475 540
rect 2205 360 2250 405
<< end >>
